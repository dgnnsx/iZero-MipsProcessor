module memoria_de_instrucoes (clk, we, addr, datain, dataout);
	input clk;										// clock
	input we;										// write enable
	input [25:0] addr;							// ram address
	input [31:0] datain;							// data in (to memory)
	
	output [31:0] dataout;						// data out (from memory)
	
	parameter RAM_SIZE = 71;					// Tamanho da memoria
	reg [31:0] ram [RAM_SIZE-1:0];			// ram cells
	
	assign dataout = ram[addr];				// use 5-bit word address
	
	always @ (posedge clk) begin
		if (we) ram[addr] <= datain;			// write ram
	end

	integer i;
	initial begin
		// ram initialization
		//for (i = 0; i < RAM_SIZE; i = i + 1)
			//ram[i] <= 0;
			ram[0] <= 32'b010110_00000000000000000000101110;		// Jump to Main
			ram[1] <= 32'b000001_11110_11110_0000000000001000; 	// addi
			ram[2] <= 32'b010010_11110_00110_1111111111111011; 	// sw
			ram[3] <= 32'b010010_11110_00111_1111111111111100; 	// sw
			ram[4] <= 32'b010000_00000_10100_0000000000000000; 	// li
			ram[5] <= 32'b010010_11110_10100_1111111111111101; 	// sw
			ram[6] <= 32'b001111_11110_01010_1111111111111100; 	// lw
			ram[7] <= 32'b000010_01010_10101_0000000000000001; 	// subi
			ram[8] <= 32'b001111_11110_01011_1111111111111101; 	// lw
			ram[9] <= 32'b000000_01011_10101_10110_00000_001110; 	// lt
			ram[10] <= 32'b010101_10110_00000_0000000000101101; 	// jf
			ram[11] <= 32'b010010_11110_01011_1111111111111111; 	// sw
			ram[12] <= 32'b000001_01011_10111_0000000000000001; 	// addi
			ram[13] <= 32'b010010_11110_10111_1111111111111110; 	// sw
			ram[14] <= 32'b001111_11110_01100_1111111111111110; 	// lw
			ram[15] <= 32'b000000_01100_01010_11000_00000_001110; 	// lt
			ram[16] <= 32'b010101_11000_00000_0000000000011101; 	// jf
			ram[17] <= 32'b001111_11110_01101_1111111111111011; 	// lw
			ram[18] <= 32'b000000_01101_01100_11001_00000_000000; 	// add
			ram[19] <= 32'b001111_11001_11001_0000000000000000; 	// lw
			ram[20] <= 32'b001111_11110_01110_1111111111111111; 	// lw
			ram[21] <= 32'b000000_01101_01110_11010_00000_000000; 	// add
			ram[22] <= 32'b001111_11010_11010_0000000000000000; 	// lw
			ram[23] <= 32'b000000_11001_11010_11011_00000_001110; 	// lt
			ram[24] <= 32'b010101_11011_00000_0000000000011010; 	// jf
			ram[25] <= 32'b010010_11110_01100_1111111111111111; 	// sw
			ram[26] <= 32'b000001_01100_11100_0000000000000001; 	// addi
			ram[27] <= 32'b010010_11110_11100_1111111111111110; 	// sw
			ram[28] <= 32'b010110_00000000000000000000001110; 	// j
			ram[29] <= 32'b001111_11110_01111_1111111111111111; 	// lw
			ram[30] <= 32'b000000_01011_01111_11101_00000_001101; 	// ne
			ram[31] <= 32'b010101_11101_00000_0000000000101010; 	// jf
			ram[32] <= 32'b000000_01101_01011_10100_00000_000000; 	// add
			ram[33] <= 32'b001111_10100_10100_0000000000000000; 	// lw
			ram[34] <= 32'b010010_11110_10100_0000000000000000; 	// sw
			ram[35] <= 32'b000000_01101_01111_10101_00000_000000; 	// add
			ram[36] <= 32'b001111_10101_10101_0000000000000000; 	// lw
			ram[37] <= 32'b000000_01101_01011_10110_00000_000000; 	// add
			ram[38] <= 32'b010010_10110_10101_0000000000000000; 	// sw
			ram[39] <= 32'b000000_01101_01111_10111_00000_000000; 	// add
			ram[40] <= 32'b001111_11110_10000_0000000000000000; 	// lw
			ram[41] <= 32'b010010_10111_10000_0000000000000000; 	// sw
			ram[42] <= 32'b000001_01011_11000_0000000000000001; 	// addi
			ram[43] <= 32'b010010_11110_11000_1111111111111101; 	// sw
			ram[44] <= 32'b010110_00000000000000000000000110; 	// j
			ram[45] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
			ram[46] <= 32'b000001_11110_11110_0000000000000101; 	// addi
			ram[47] <= 32'b010001_11110_01010_1111111111111100; 	// la
			ram[48] <= 32'b010000_00000_10100_0000000000001001; 	// li
			ram[49] <= 32'b010010_01010_10100_0000000000000000; 	// sw
			ram[50] <= 32'b010000_00000_10101_0000000000000110; 	// li
			ram[51] <= 32'b010010_01010_10101_0000000000000001; 	// sw
			ram[52] <= 32'b010000_00000_10110_0000000000001000; 	// li
			ram[53] <= 32'b010010_01010_10110_0000000000000010; 	// sw
			ram[54] <= 32'b010000_00000_10111_0000000000000111; 	// li
			ram[55] <= 32'b010010_01010_10111_0000000000000011; 	// sw
			ram[56] <= 32'b010001_11110_00110_1111111111111100; 	// la
			ram[57] <= 32'b010000_00000_00111_0000000000000100; 	// li
			ram[58] <= 32'b010111_00000000000000000000000001; 	// jal
			ram[59] <= 32'b001110_00001_01011_0000000000000000; 	// mov
			ram[60] <= 32'b000010_11110_11110_0000000000001000; 	// subi
			ram[61] <= 32'b010011_00000_11000_0000000000000000; 	// in
			ram[62] <= 32'b010010_11110_11000_0000000000000000; 	// sw
			ram[63] <= 32'b010001_11110_01100_1111111111111100; 	// la
			ram[64] <= 32'b001111_11110_01101_0000000000000000; 	// lw
			ram[65] <= 32'b000000_01100_01101_11001_00000_000000; 	// add
			ram[66] <= 32'b001111_11001_11001_0000000000000000; 	// lw
			ram[67] <= 32'b001110_11001_00110_0000000000000000; 	// mov
			ram[68] <= 32'b010000_00000_00111_0000000000000010; 	// li
			ram[69] <= 32'b010100_00000_00110_0000000000000010; 	// out
			ram[70] <= 32'b011000_00000000000000000000000000; 	// halt
	end
endmodule
