module bios(pc, instrucao);
	// Entrada
	input [25:0] pc;										// PC Atual
	
	// Saida
	output [31:0] instrucao;							// Proxima instrucao a ser executada
	
	localparam BIOS_SIZE = 52;							// Tamanho da bios
	wire [31:0] bios [BIOS_SIZE-1:0];				// Memoria da bios
	
	assign bios[0] = 32'b010110_00000000000000000000100100;		// Jump to Main
	assign bios[1] = 32'b000001_11110_11110_0000000000000010; 	// addi
	assign bios[2] = 32'b011101_00000000000000000000000000; 	// ckhd
	assign bios[3] = 32'b011110_00000000000000000000000000; 	// ckim
	assign bios[4] = 32'b011111_00000000000000000000000000; 	// ckdm
	assign bios[5] = 32'b000000_11111_00000_00000_00000_010010; 	// jr
	assign bios[6] = 32'b000001_11110_11110_0000000000000101; 	// addi
	assign bios[7] = 32'b010000_00000_10100_0000000000011000; 	// li
	assign bios[8] = 32'b010010_11110_10100_0000000000000000; 	// sw
	assign bios[9] = 32'b010000_00000_10101_0000000000000000; 	// li
	assign bios[10] = 32'b010010_11110_10101_1111111111111111; 	// sw
	assign bios[11] = 32'b001111_11110_01010_1111111111111111; 	// lw
	assign bios[12] = 32'b001110_01010_00110_0000000000000000; 	// mov
	assign bios[13] = 32'b011001_00110_10110_0000000000000000; 	// ldk
	assign bios[14] = 32'b010010_11110_10110_1111111111111110; 	// sw
	assign bios[15] = 32'b001111_11110_01011_1111111111111110; 	// lw
	assign bios[16] = 32'b001101_01011_10111_0000000000011010; 	// srli
	assign bios[17] = 32'b001111_11110_01100_0000000000000000; 	// lw
	assign bios[18] = 32'b000000_10111_01100_11000_00000_001101; 	// ne
	assign bios[19] = 32'b010101_11000_00000_0000000000011111; 	// jf
	assign bios[20] = 32'b001110_01011_00110_0000000000000000; 	// mov
	assign bios[21] = 32'b001110_01010_00111_0000000000000000; 	// mov
	assign bios[22] = 32'b011100_00111_00110_0000000000000000; 	// sim
	assign bios[23] = 32'b000001_01010_11001_0000000000000001; 	// addi
	assign bios[24] = 32'b010010_11110_11001_1111111111111111; 	// sw
	assign bios[25] = 32'b001111_11110_01010_1111111111111111; 	// lw
	assign bios[26] = 32'b001110_01010_00110_0000000000000000; 	// mov
	assign bios[27] = 32'b011001_00110_11010_0000000000000000; 	// ldk
	assign bios[28] = 32'b010010_11110_11010_1111111111111110; 	// sw
	assign bios[29] = 32'b001111_11110_01011_1111111111111110; 	// lw
	assign bios[30] = 32'b010110_00000000000000000000001111; 	// j
	assign bios[31] = 32'b001110_01011_00110_0000000000000000; 	// mov
	assign bios[32] = 32'b001110_01010_00111_0000000000000000; 	// mov
	assign bios[33] = 32'b011100_00111_00110_0000000000000000; 	// sim
	assign bios[34] = 32'b001110_01010_00001_0000000000000000; 	// mov
	assign bios[35] = 32'b000000_11111_00000_00000_00000_010010; 	// jr
	assign bios[36] = 32'b000001_11110_11110_0000000000000011; 	// addi
	assign bios[37] = 32'b010111_00000000000000000000000110; 	// jal
	assign bios[38] = 32'b001110_00001_01010_0000000000000000; 	// mov
	assign bios[39] = 32'b000010_11110_11110_0000000000000101; 	// subi
	assign bios[40] = 32'b010010_11110_01010_0000000000000000; 	// sw
	assign bios[41] = 32'b010000_00000_10100_0000000000000000; 	// li
	assign bios[42] = 32'b010010_11110_10100_1111111111111110; 	// sw
	assign bios[43] = 32'b001111_11110_01011_0000000000000000; 	// lw
	assign bios[44] = 32'b010010_11110_01011_1111111111111111; 	// sw
	assign bios[45] = 32'b001111_11110_01100_1111111111111110; 	// lw
	assign bios[46] = 32'b001110_01100_00110_0000000000000000; 	// mov
	assign bios[47] = 32'b010000_00000_00111_0000000000000000; 	// li
	assign bios[48] = 32'b100000_00111_00110_0000000000000000; 	// mmuLower
	assign bios[49] = 32'b011000_00000000000000000000000000; 	// halt

	assign instrucao = bios[pc];
endmodule
