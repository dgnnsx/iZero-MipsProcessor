library verilog;
use verilog.vl_types.all;
entity memoria_de_dados_vlg_vec_tst is
end memoria_de_dados_vlg_vec_tst;
