module disco_rigido (clk, we, addr, datain, dataout);
	input clk;										// clock
	input we;										// write enable
	input [31:0] addr;							// disk address
	input [31:0] datain;							// data in (to disk)
	
	output reg [31:0] dataout;					// data out (from disk)
	
	localparam DISK_SIZE = 2048;				// Tamanho do disco
	reg [31:0] disk [DISK_SIZE-1:0];			// disk cells
	
	always @ (posedge clk) begin
		if (we) disk[addr] <= datain;			// write disk
	end
	
	always @ (negedge clk) begin
		dataout <= disk[addr];
	end

	initial begin
		// SISTEMA OPERACIONAL

disk[0] <= 32'b111100_00000000000000001101111010;		// Jump to Main
disk[1] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[2] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[3] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[4] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[5] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[6] <= 32'b010110_00001_10000_0000000000000000; 	// ldk
disk[7] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[8] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[9] <= 32'b001101_00101_10001_0000000000011010; 	// srli
disk[10] <= 32'b001111_11101_00110_0000000011111001; 	// lw
disk[11] <= 32'b000000_10001_00110_10010_00000_001101; 	// ne
disk[12] <= 32'b010101_10010_00000_0000000000010110; 	// jf
disk[13] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[14] <= 32'b000001_00111_10011_0000000000000001; 	// addi
disk[15] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[16] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[17] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[18] <= 32'b010110_00001_10100_0000000000000000; 	// ldk
disk[19] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[20] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[21] <= 32'b111100_00000000000000000000001000; 	// j
disk[22] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[23] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[24] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[25] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[26] <= 32'b010010_11110_00001_1111111111111111; 	// sw
disk[27] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[28] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[29] <= 32'b000000_00101_10000_01111_00000_001100; 	// eq
disk[30] <= 32'b010101_01111_00000_0000000000100010; 	// jf
disk[31] <= 32'b010000_00000_10001_0000000000000001; 	// li
disk[32] <= 32'b001110_10001_11001_0000000000000000; 	// mov
disk[33] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[34] <= 32'b010000_00000_10010_0000000000000001; 	// li
disk[35] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[36] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[37] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[38] <= 32'b000000_00101_10100_10011_00000_010000; 	// gt
disk[39] <= 32'b010101_10011_00000_0000000000110000; 	// jf
disk[40] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[41] <= 32'b000011_00110_10101_0000000000000010; 	// muli
disk[42] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[43] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[44] <= 32'b000010_00101_10110_0000000000000001; 	// subi
disk[45] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[46] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[47] <= 32'b111100_00000000000000000000100100; 	// j
disk[48] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[49] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[50] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[51] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[52] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[53] <= 32'b010000_00000_00010_0000000000000000; 	// li
disk[54] <= 32'b010100_00000_00001_0000000000000000; 	// out
disk[55] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[56] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[57] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[58] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[59] <= 32'b010000_00000_00010_0000000000000010; 	// li
disk[60] <= 32'b010100_00000_00001_0000000000000010; 	// out
disk[61] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[62] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[63] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[64] <= 32'b010010_11101_01111_0000000011001010; 	// sw
disk[65] <= 32'b010000_00000_10000_0000000000000001; 	// li
disk[66] <= 32'b010010_11101_10000_0000000011001011; 	// sw
disk[67] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[68] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[69] <= 32'b010000_00000_01111_0000000000000001; 	// li
disk[70] <= 32'b010010_11101_01111_0000000000000000; 	// sw
disk[71] <= 32'b010000_00000_10000_0000000000000010; 	// li
disk[72] <= 32'b010010_11101_10000_0000000000000001; 	// sw
disk[73] <= 32'b010000_00000_10001_0000000000000011; 	// li
disk[74] <= 32'b010010_11101_10001_0000000000000010; 	// sw
disk[75] <= 32'b010000_00000_10010_0000000110010100; 	// li
disk[76] <= 32'b010010_11101_10010_0000000000000011; 	// sw
disk[77] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[78] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[79] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[80] <= 32'b010000_00000_10101_0000000000001010; 	// li
disk[81] <= 32'b000000_00101_10101_10100_00000_001110; 	// lt
disk[82] <= 32'b010101_10100_00000_0000000001101111; 	// jf
disk[83] <= 32'b010001_11101_00110_0000000000000100; 	// la
disk[84] <= 32'b000000_00110_00101_10110_00000_000000; 	// add
disk[85] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[86] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[87] <= 32'b010001_11101_00111_0000000000001110; 	// la
disk[88] <= 32'b000000_00111_00101_11000_00000_000000; 	// add
disk[89] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[90] <= 32'b010010_11000_01111_0000000000000000; 	// sw
disk[91] <= 32'b010001_11101_01000_0000000000011000; 	// la
disk[92] <= 32'b000000_01000_00101_10000_00000_000000; 	// add
disk[93] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[94] <= 32'b010010_10000_10001_0000000000000000; 	// sw
disk[95] <= 32'b010001_11101_01001_0000000000100010; 	// la
disk[96] <= 32'b000000_01001_00101_10010_00000_000000; 	// add
disk[97] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[98] <= 32'b010010_10010_10011_0000000000000000; 	// sw
disk[99] <= 32'b010001_11101_01010_0000000000101100; 	// la
disk[100] <= 32'b000000_01010_00101_10100_00000_000000; 	// add
disk[101] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[102] <= 32'b010010_10100_10101_0000000000000000; 	// sw
disk[103] <= 32'b010001_11101_01011_0000000000110110; 	// la
disk[104] <= 32'b000000_01011_00101_10110_00000_000000; 	// add
disk[105] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[106] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[107] <= 32'b000001_00101_11000_0000000000000001; 	// addi
disk[108] <= 32'b010010_11110_11000_0000000000000000; 	// sw
disk[109] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[110] <= 32'b111100_00000000000000000001001111; 	// j
disk[111] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[112] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[113] <= 32'b010000_00000_01111_0000000000100000; 	// li
disk[114] <= 32'b010010_11101_01111_0000000010000010; 	// sw
disk[115] <= 32'b010000_00000_10000_0000000001000000; 	// li
disk[116] <= 32'b010010_11101_10000_0000000010000011; 	// sw
disk[117] <= 32'b010000_00000_10001_0000000001100100; 	// li
disk[118] <= 32'b010010_11101_10001_0000000010000100; 	// sw
disk[119] <= 32'b010000_00000_10010_0000000000001010; 	// li
disk[120] <= 32'b010010_11101_10010_0000000010000101; 	// sw
disk[121] <= 32'b010000_00000_10011_0000001111100111; 	// li
disk[122] <= 32'b010010_11101_10011_0000000001000000; 	// sw
disk[123] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[124] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[125] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[126] <= 32'b010010_11101_01111_0000000011111010; 	// sw
disk[127] <= 32'b010000_00000_10000_0000000000000001; 	// li
disk[128] <= 32'b010010_11101_10000_0000000011111011; 	// sw
disk[129] <= 32'b010000_00000_10001_0000000000000010; 	// li
disk[130] <= 32'b010010_11101_10001_0000000011111100; 	// sw
disk[131] <= 32'b010000_00000_10010_0000000000000011; 	// li
disk[132] <= 32'b010010_11101_10010_0000000011111101; 	// sw
disk[133] <= 32'b010000_00000_10011_0000000000000100; 	// li
disk[134] <= 32'b010010_11101_10011_0000000011111110; 	// sw
disk[135] <= 32'b010000_00000_10100_0000000000000101; 	// li
disk[136] <= 32'b010010_11101_10100_0000000011111111; 	// sw
disk[137] <= 32'b010000_00000_10101_0000000000000110; 	// li
disk[138] <= 32'b010010_11101_10101_0000000100000000; 	// sw
disk[139] <= 32'b010000_00000_10110_0000000000011110; 	// li
disk[140] <= 32'b010010_11101_10110_0000000100000001; 	// sw
disk[141] <= 32'b001111_11101_00101_0000000011111010; 	// lw
disk[142] <= 32'b010010_11101_00101_0000000100000010; 	// sw
disk[143] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[144] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[145] <= 32'b010000_00000_01111_0000011111111111; 	// li
disk[146] <= 32'b010010_11101_01111_0000000010000111; 	// sw
disk[147] <= 32'b010000_00000_10000_0000000000011111; 	// li
disk[148] <= 32'b010010_11101_10000_0000000011110111; 	// sw
disk[149] <= 32'b010000_00000_10001_0000000000111101; 	// li
disk[150] <= 32'b010010_11101_10001_0000000011111000; 	// sw
disk[151] <= 32'b010000_00000_10010_0000000000111111; 	// li
disk[152] <= 32'b010010_11101_10010_0000000011111001; 	// sw
disk[153] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[154] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[155] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[156] <= 32'b010010_11110_01111_1111111111111110; 	// sw
disk[157] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[158] <= 32'b001111_11101_00110_0000000010000011; 	// lw
disk[159] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[160] <= 32'b010101_10000_00000_0000000010101101; 	// jf
disk[161] <= 32'b010001_11101_00111_0000000001000010; 	// la
disk[162] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[163] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[164] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[165] <= 32'b010001_11101_01000_0000000010001010; 	// la
disk[166] <= 32'b000000_01000_00101_10011_00000_000000; 	// add
disk[167] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[168] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[169] <= 32'b000001_00101_10101_0000000000000001; 	// addi
disk[170] <= 32'b010010_11110_10101_1111111111111110; 	// sw
disk[171] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[172] <= 32'b111100_00000000000000000010011101; 	// j
disk[173] <= 32'b010010_11110_11111_1111111111111101; 	// sw
disk[174] <= 32'b111110_00000000000000000000000001; 	// jal
disk[175] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[176] <= 32'b001111_11110_11111_1111111111111101; 	// lw
disk[177] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[178] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[179] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[180] <= 32'b000001_00110_10110_0000000000000001; 	// addi
disk[181] <= 32'b010010_11101_10110_0000000010000110; 	// sw
disk[182] <= 32'b001111_11101_00111_0000000010000010; 	// lw
disk[183] <= 32'b000000_00110_00111_10111_00000_000011; 	// div
disk[184] <= 32'b010010_11110_10111_1111111111111111; 	// sw
disk[185] <= 32'b000000_00110_00111_11000_00000_000100; 	// mod
disk[186] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[187] <= 32'b000000_11000_10000_01111_00000_010000; 	// gt
disk[188] <= 32'b010101_01111_00000_0000000011000001; 	// jf
disk[189] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[190] <= 32'b000001_01000_10001_0000000000000001; 	// addi
disk[191] <= 32'b010010_11110_10001_1111111111111111; 	// sw
disk[192] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[193] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[194] <= 32'b010010_11110_10010_1111111111111110; 	// sw
disk[195] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[196] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[197] <= 32'b000000_00101_00110_10011_00000_001110; 	// lt
disk[198] <= 32'b010101_10011_00000_0000000011001111; 	// jf
disk[199] <= 32'b010001_11101_00111_0000000001000010; 	// la
disk[200] <= 32'b000000_00111_00101_10100_00000_000000; 	// add
disk[201] <= 32'b010000_00000_10101_0000000000000001; 	// li
disk[202] <= 32'b010010_10100_10101_0000000000000000; 	// sw
disk[203] <= 32'b000001_00101_10110_0000000000000001; 	// addi
disk[204] <= 32'b010010_11110_10110_1111111111111110; 	// sw
disk[205] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[206] <= 32'b111100_00000000000000000011000011; 	// j
disk[207] <= 32'b001110_11110_10111_0000000000000000; 	// mov
disk[208] <= 32'b001111_11101_00101_0000000010000010; 	// lw
disk[209] <= 32'b000000_10111_00101_11000_00000_000011; 	// div
disk[210] <= 32'b010010_11110_11000_1111111111111111; 	// sw
disk[211] <= 32'b001110_11110_01111_0000000000000000; 	// mov
disk[212] <= 32'b000000_01111_00101_10000_00000_000100; 	// mod
disk[213] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[214] <= 32'b000000_10000_10010_10001_00000_010000; 	// gt
disk[215] <= 32'b010101_10001_00000_0000000011011100; 	// jf
disk[216] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[217] <= 32'b000001_00110_10011_0000000000000001; 	// addi
disk[218] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[219] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[220] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[221] <= 32'b010010_11110_10100_1111111111111110; 	// sw
disk[222] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[223] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[224] <= 32'b000000_00101_00110_10101_00000_001110; 	// lt
disk[225] <= 32'b010101_10101_00000_0000000011101010; 	// jf
disk[226] <= 32'b010001_11101_00111_0000000010001010; 	// la
disk[227] <= 32'b000000_00111_00101_10110_00000_000000; 	// add
disk[228] <= 32'b010000_00000_10111_0000000000000001; 	// li
disk[229] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[230] <= 32'b000001_00101_11000_0000000000000001; 	// addi
disk[231] <= 32'b010010_11110_11000_1111111111111110; 	// sw
disk[232] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[233] <= 32'b111100_00000000000000000011011110; 	// j
disk[234] <= 32'b001111_11101_00101_0000000010000011; 	// lw
disk[235] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[236] <= 32'b010001_11101_00110_0000000010001010; 	// la
disk[237] <= 32'b000000_00110_01111_10000_00000_000000; 	// add
disk[238] <= 32'b010000_00000_10001_0000000000000001; 	// li
disk[239] <= 32'b010010_10000_10001_0000000000000000; 	// sw
disk[240] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[241] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[242] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[243] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[244] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[245] <= 32'b001111_11101_00110_0000000010000101; 	// lw
disk[246] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[247] <= 32'b010101_10000_00000_0000000100001100; 	// jf
disk[248] <= 32'b010001_11101_00111_0000000011001111; 	// la
disk[249] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[250] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[251] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[252] <= 32'b010001_11101_01000_0000000011011001; 	// la
disk[253] <= 32'b000000_01000_00101_10011_00000_000000; 	// add
disk[254] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[255] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[256] <= 32'b010001_11101_01001_0000000011100011; 	// la
disk[257] <= 32'b000000_01001_00101_10101_00000_000000; 	// add
disk[258] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[259] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[260] <= 32'b010001_11101_01010_0000000011101101; 	// la
disk[261] <= 32'b000000_01010_00101_10111_00000_000000; 	// add
disk[262] <= 32'b010000_00000_11000_0000000000000000; 	// li
disk[263] <= 32'b010010_10111_11000_0000000000000000; 	// sw
disk[264] <= 32'b000001_00101_01111_0000000000000001; 	// addi
disk[265] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[266] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[267] <= 32'b111100_00000000000000000011110100; 	// j
disk[268] <= 32'b001111_11101_00101_0000000010000110; 	// lw
disk[269] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[270] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[271] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[272] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[273] <= 32'b001111_11101_00110_0000000010000111; 	// lw
disk[274] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[275] <= 32'b010101_10001_00000_0000000100101100; 	// jf
disk[276] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[277] <= 32'b010110_00001_10010_0000000000000000; 	// ldk
disk[278] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[279] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[280] <= 32'b001101_00111_10011_0000000000011010; 	// srli
disk[281] <= 32'b001111_11101_01000_0000000011111000; 	// lw
disk[282] <= 32'b000000_10011_01000_10100_00000_001100; 	// eq
disk[283] <= 32'b010101_10100_00000_0000000100100111; 	// jf
disk[284] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[285] <= 32'b000001_01001_10101_0000000000000001; 	// addi
disk[286] <= 32'b010001_11101_01010_0000000011001111; 	// la
disk[287] <= 32'b000000_01010_01001_10110_00000_000000; 	// add
disk[288] <= 32'b010010_10110_10101_0000000000000000; 	// sw
disk[289] <= 32'b010001_11101_01011_0000000011011001; 	// la
disk[290] <= 32'b000000_01011_01001_10111_00000_000000; 	// add
disk[291] <= 32'b010010_10111_00101_0000000000000000; 	// sw
disk[292] <= 32'b000001_01001_11000_0000000000000001; 	// addi
disk[293] <= 32'b010010_11110_11000_1111111111111111; 	// sw
disk[294] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[295] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[296] <= 32'b000001_00101_01111_0000000000000001; 	// addi
disk[297] <= 32'b010010_11110_01111_1111111111111110; 	// sw
disk[298] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[299] <= 32'b111100_00000000000000000100010000; 	// j
disk[300] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[301] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[302] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[303] <= 32'b111110_00000000000000000001000100; 	// jal
disk[304] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[305] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[306] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[307] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[308] <= 32'b111110_00000000000000000001110000; 	// jal
disk[309] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[310] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[311] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[312] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[313] <= 32'b111110_00000000000000000001111100; 	// jal
disk[314] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[315] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[316] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[317] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[318] <= 32'b111110_00000000000000000010010000; 	// jal
disk[319] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[320] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[321] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[322] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[323] <= 32'b111110_00000000000000000010011010; 	// jal
disk[324] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[325] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[326] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[327] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[328] <= 32'b111110_00000000000000000011110001; 	// jal
disk[329] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[330] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[331] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[332] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[333] <= 32'b000001_11110_11110_0000000000000110; 	// addi
disk[334] <= 32'b010010_11110_00001_1111111111111101; 	// sw
disk[335] <= 32'b001111_11110_00101_1111111111111101; 	// lw
disk[336] <= 32'b001111_11101_00110_0000000010000010; 	// lw
disk[337] <= 32'b000000_00101_00110_01111_00000_000011; 	// div
disk[338] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[339] <= 32'b000000_00101_00110_10000_00000_000100; 	// mod
disk[340] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[341] <= 32'b000000_10000_10010_10001_00000_010000; 	// gt
disk[342] <= 32'b010101_10001_00000_0000000101011011; 	// jf
disk[343] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[344] <= 32'b000001_00111_10011_0000000000000001; 	// addi
disk[345] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[346] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[347] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[348] <= 32'b010010_11110_10100_1111111111111110; 	// sw
disk[349] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[350] <= 32'b001111_11101_00110_0000000010000011; 	// lw
disk[351] <= 32'b000000_00101_00110_10101_00000_001110; 	// lt
disk[352] <= 32'b010101_10101_00000_0000000110000000; 	// jf
disk[353] <= 32'b010001_11101_00111_0000000001000010; 	// la
disk[354] <= 32'b000000_00111_00101_10110_00000_000000; 	// add
disk[355] <= 32'b001111_10110_10110_0000000000000000; 	// lw
disk[356] <= 32'b010000_00000_11000_0000000000000000; 	// li
disk[357] <= 32'b000000_10110_11000_10111_00000_001100; 	// eq
disk[358] <= 32'b010101_10111_00000_0000000101111011; 	// jf
disk[359] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[360] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[361] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[362] <= 32'b000000_00101_10000_01111_00000_010000; 	// gt
disk[363] <= 32'b010101_01111_00000_0000000101111000; 	// jf
disk[364] <= 32'b010001_11101_00110_0000000001000010; 	// la
disk[365] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[366] <= 32'b000000_00110_00111_10001_00000_000000; 	// add
disk[367] <= 32'b010000_00000_10010_0000000000000001; 	// li
disk[368] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[369] <= 32'b000010_00101_10011_0000000000000001; 	// subi
disk[370] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[371] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[372] <= 32'b000001_00111_10100_0000000000000001; 	// addi
disk[373] <= 32'b010010_11110_10100_1111111111111110; 	// sw
disk[374] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[375] <= 32'b111100_00000000000000000101101000; 	// j
disk[376] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[377] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[378] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[379] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[380] <= 32'b000001_00101_10101_0000000000000001; 	// addi
disk[381] <= 32'b010010_11110_10101_1111111111111110; 	// sw
disk[382] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[383] <= 32'b111100_00000000000000000101011101; 	// j
disk[384] <= 32'b001111_11101_00101_0000000010000100; 	// lw
disk[385] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[386] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[387] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[388] <= 32'b010001_11101_00101_0000000000101100; 	// la
disk[389] <= 32'b001111_11101_00110_0000000001000001; 	// lw
disk[390] <= 32'b000000_00101_00110_01111_00000_000000; 	// add
disk[391] <= 32'b001111_01111_01111_0000000000000000; 	// lw
disk[392] <= 32'b001111_11101_00111_0000000010000010; 	// lw
disk[393] <= 32'b000000_01111_00111_10000_00000_000011; 	// div
disk[394] <= 32'b000001_10000_10001_0000000000000001; 	// addi
disk[395] <= 32'b010010_11110_10001_1111111111111111; 	// sw
disk[396] <= 32'b000000_00101_00110_10010_00000_000000; 	// add
disk[397] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[398] <= 32'b000000_10010_00111_10011_00000_000100; 	// mod
disk[399] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[400] <= 32'b000000_10011_10101_10100_00000_010000; 	// gt
disk[401] <= 32'b010101_10100_00000_0000000110010110; 	// jf
disk[402] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[403] <= 32'b000001_01000_10110_0000000000000001; 	// addi
disk[404] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[405] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[406] <= 32'b001111_11101_00101_0000000010000011; 	// lw
disk[407] <= 32'b000010_00101_10111_0000000000000001; 	// subi
disk[408] <= 32'b010010_11110_10111_1111111111111110; 	// sw
disk[409] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[410] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[411] <= 32'b000000_00101_01111_11000_00000_010000; 	// gt
disk[412] <= 32'b010101_11000_00000_0000000110111100; 	// jf
disk[413] <= 32'b010001_11101_00110_0000000010001010; 	// la
disk[414] <= 32'b000000_00110_00101_10000_00000_000000; 	// add
disk[415] <= 32'b001111_10000_10000_0000000000000000; 	// lw
disk[416] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[417] <= 32'b000000_10000_10010_10001_00000_001100; 	// eq
disk[418] <= 32'b010101_10001_00000_0000000110110111; 	// jf
disk[419] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[420] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[421] <= 32'b000000_00101_10100_10011_00000_010000; 	// gt
disk[422] <= 32'b010101_10011_00000_0000000110110100; 	// jf
disk[423] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[424] <= 32'b010010_11110_00110_0000000000000000; 	// sw
disk[425] <= 32'b010001_11101_00111_0000000010001010; 	// la
disk[426] <= 32'b000000_00111_00110_10101_00000_000000; 	// add
disk[427] <= 32'b010000_00000_10110_0000000000000001; 	// li
disk[428] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[429] <= 32'b000010_00101_10111_0000000000000001; 	// subi
disk[430] <= 32'b010010_11110_10111_1111111111111111; 	// sw
disk[431] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[432] <= 32'b000010_00110_11000_0000000000000001; 	// subi
disk[433] <= 32'b010010_11110_11000_1111111111111110; 	// sw
disk[434] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[435] <= 32'b111100_00000000000000000110100011; 	// j
disk[436] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[437] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[438] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[439] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[440] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[441] <= 32'b010010_11110_01111_1111111111111110; 	// sw
disk[442] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[443] <= 32'b111100_00000000000000000110011001; 	// j
disk[444] <= 32'b001111_11101_00101_0000000010000100; 	// lw
disk[445] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[446] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[447] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[448] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[449] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[450] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[451] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[452] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[453] <= 32'b001111_11101_00110_0000000010000101; 	// lw
disk[454] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[455] <= 32'b010101_10001_00000_0000000111011101; 	// jf
disk[456] <= 32'b010001_11101_00111_0000000011100011; 	// la
disk[457] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
disk[458] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[459] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[460] <= 32'b000000_10010_10100_10011_00000_001101; 	// ne
disk[461] <= 32'b010101_10011_00000_0000000111011000; 	// jf
disk[462] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[463] <= 32'b010010_11110_11111_1111111111111110; 	// sw
disk[464] <= 32'b111110_00000000000000000000011001; 	// jal
disk[465] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[466] <= 32'b001111_11110_11111_1111111111111110; 	// lw
disk[467] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[468] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[469] <= 32'b000000_00110_00101_10101_00000_000000; 	// add
disk[470] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[471] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[472] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[473] <= 32'b000001_00101_10110_0000000000000001; 	// addi
disk[474] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[475] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[476] <= 32'b111100_00000000000000000111000100; 	// j
disk[477] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[478] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[479] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[480] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[481] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[482] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[483] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[484] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[485] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[486] <= 32'b001111_11101_00110_0000000010000101; 	// lw
disk[487] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[488] <= 32'b010101_10001_00000_0000000111111110; 	// jf
disk[489] <= 32'b010001_11101_00111_0000000011001111; 	// la
disk[490] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
disk[491] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[492] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[493] <= 32'b000000_10010_10100_10011_00000_001101; 	// ne
disk[494] <= 32'b010101_10011_00000_0000000111111001; 	// jf
disk[495] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[496] <= 32'b010010_11110_11111_1111111111111110; 	// sw
disk[497] <= 32'b111110_00000000000000000000011001; 	// jal
disk[498] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[499] <= 32'b001111_11110_11111_1111111111111110; 	// lw
disk[500] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[501] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[502] <= 32'b000000_00110_00101_10101_00000_000000; 	// add
disk[503] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[504] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[505] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[506] <= 32'b000001_00101_10110_0000000000000001; 	// addi
disk[507] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[508] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[509] <= 32'b111100_00000000000000000111100101; 	// j
disk[510] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[511] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[512] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[513] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[514] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[515] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[516] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[517] <= 32'b001111_11101_00110_0000000010000101; 	// lw
disk[518] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[519] <= 32'b010101_10000_00000_0000001000010101; 	// jf
disk[520] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[521] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[522] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[523] <= 32'b001111_11101_01000_0000000000000010; 	// lw
disk[524] <= 32'b000000_10001_01000_10010_00000_001100; 	// eq
disk[525] <= 32'b010101_10010_00000_0000001000010000; 	// jf
disk[526] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[527] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[528] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[529] <= 32'b000001_00101_10011_0000000000000001; 	// addi
disk[530] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[531] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[532] <= 32'b111100_00000000000000001000000100; 	// j
disk[533] <= 32'b001111_11101_00101_0000000000000011; 	// lw
disk[534] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[535] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[536] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[537] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[538] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[539] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[540] <= 32'b001111_11101_00110_0000000010000101; 	// lw
disk[541] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[542] <= 32'b010101_10000_00000_0000001000101100; 	// jf
disk[543] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[544] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[545] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[546] <= 32'b001111_11101_01000_0000000000000001; 	// lw
disk[547] <= 32'b000000_10001_01000_10010_00000_001100; 	// eq
disk[548] <= 32'b010101_10010_00000_0000001000100111; 	// jf
disk[549] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[550] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[551] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[552] <= 32'b000001_00101_10011_0000000000000001; 	// addi
disk[553] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[554] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[555] <= 32'b111100_00000000000000001000011011; 	// j
disk[556] <= 32'b001111_11101_00101_0000000000000011; 	// lw
disk[557] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[558] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[559] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[560] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[561] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[562] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[563] <= 32'b001111_11101_00110_0000000010000101; 	// lw
disk[564] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[565] <= 32'b010101_10000_00000_0000001001000101; 	// jf
disk[566] <= 32'b010001_11101_00111_0000000011100011; 	// la
disk[567] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[568] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[569] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[570] <= 32'b000000_10001_10011_10010_00000_001101; 	// ne
disk[571] <= 32'b010101_10010_00000_0000001001000000; 	// jf
disk[572] <= 32'b010001_11101_01000_0000000000000100; 	// la
disk[573] <= 32'b000000_01000_00101_10100_00000_000000; 	// add
disk[574] <= 32'b001111_11101_01001_0000000000000001; 	// lw
disk[575] <= 32'b010010_10100_01001_0000000000000000; 	// sw
disk[576] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[577] <= 32'b000001_00101_10101_0000000000000001; 	// addi
disk[578] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[579] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[580] <= 32'b111100_00000000000000001000110010; 	// j
disk[581] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[582] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[583] <= 32'b010010_11110_00001_1111111111111110; 	// sw
disk[584] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[585] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[586] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[587] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[588] <= 32'b010110_00001_01111_0000000000000000; 	// ldk
disk[589] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[590] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[591] <= 32'b001101_00101_10000_0000000000011010; 	// srli
disk[592] <= 32'b001111_11101_00110_0000000011110111; 	// lw
disk[593] <= 32'b000000_10000_00110_10001_00000_001101; 	// ne
disk[594] <= 32'b010101_10001_00000_0000001001011100; 	// jf
disk[595] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[596] <= 32'b000001_00111_10010_0000000000000001; 	// addi
disk[597] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[598] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[599] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[600] <= 32'b010110_00001_10011_0000000000000000; 	// ldk
disk[601] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[602] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[603] <= 32'b111100_00000000000000001001001110; 	// j
disk[604] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[605] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[606] <= 32'b000000_00101_00110_10100_00000_000001; 	// sub
disk[607] <= 32'b001110_10100_11001_0000000000000000; 	// mov
disk[608] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[609] <= 32'b000001_11110_11110_0000000000001010; 	// addi
disk[610] <= 32'b010010_11110_00001_1111111111111001; 	// sw
disk[611] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[612] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[613] <= 32'b010010_11110_01111_1111111111111001; 	// sw
disk[614] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[615] <= 32'b010001_11101_00110_0000000011011001; 	// la
disk[616] <= 32'b000000_00110_00101_10000_00000_000000; 	// add
disk[617] <= 32'b001111_10000_10000_0000000000000000; 	// lw
disk[618] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[619] <= 32'b010001_11101_00111_0000000011001111; 	// la
disk[620] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[621] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[622] <= 32'b010010_11110_10001_0000000000000000; 	// sw
disk[623] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[624] <= 32'b010010_11110_01000_1111111111111010; 	// sw
disk[625] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[626] <= 32'b010010_11110_11111_1111111111111000; 	// sw
disk[627] <= 32'b111110_00000000000000001001000110; 	// jal
disk[628] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[629] <= 32'b001111_11110_11111_1111111111111000; 	// lw
disk[630] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[631] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[632] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[633] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[634] <= 32'b010010_11110_11111_1111111111111000; 	// sw
disk[635] <= 32'b111110_00000000000000000101001101; 	// jal
disk[636] <= 32'b000010_11110_11110_0000000000000110; 	// subi
disk[637] <= 32'b001111_11110_11111_1111111111111000; 	// lw
disk[638] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[639] <= 32'b010010_11110_00101_1111111111111101; 	// sw
disk[640] <= 32'b001111_11101_00110_0000000010000010; 	// lw
disk[641] <= 32'b001111_11110_00111_1111111111111101; 	// lw
disk[642] <= 32'b000000_00110_00111_10010_00000_000010; 	// mul
disk[643] <= 32'b010010_11110_10010_1111111111111011; 	// sw
disk[644] <= 32'b001111_11110_01000_1111111111111010; 	// lw
disk[645] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[646] <= 32'b010110_00001_10011_0000000000000000; 	// ldk
disk[647] <= 32'b010010_11110_10011_1111111111111100; 	// sw
disk[648] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[649] <= 32'b001101_00101_10100_0000000000011010; 	// srli
disk[650] <= 32'b001111_11101_00110_0000000011110111; 	// lw
disk[651] <= 32'b000000_10100_00110_10101_00000_001101; 	// ne
disk[652] <= 32'b010101_10101_00000_0000001010011101; 	// jf
disk[653] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[654] <= 32'b001111_11110_00111_1111111111111011; 	// lw
disk[655] <= 32'b001110_00111_00010_0000000000000000; 	// mov
disk[656] <= 32'b011001_00010_00001_0000000000000000; 	// sim
disk[657] <= 32'b001111_11110_01000_1111111111111010; 	// lw
disk[658] <= 32'b000001_01000_10110_0000000000000001; 	// addi
disk[659] <= 32'b010010_11110_10110_1111111111111010; 	// sw
disk[660] <= 32'b001111_11110_01000_1111111111111010; 	// lw
disk[661] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[662] <= 32'b010110_00001_10111_0000000000000000; 	// ldk
disk[663] <= 32'b010010_11110_10111_1111111111111100; 	// sw
disk[664] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[665] <= 32'b000001_00111_11000_0000000000000001; 	// addi
disk[666] <= 32'b010010_11110_11000_1111111111111011; 	// sw
disk[667] <= 32'b001111_11110_00111_1111111111111011; 	// lw
disk[668] <= 32'b111100_00000000000000001010001000; 	// j
disk[669] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[670] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[671] <= 32'b001111_11110_00110_1111111111111011; 	// lw
disk[672] <= 32'b001110_00110_00010_0000000000000000; 	// mov
disk[673] <= 32'b011001_00010_00001_0000000000000000; 	// sim
disk[674] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[675] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[676] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
disk[677] <= 32'b001111_11101_01000_0000000010000010; 	// lw
disk[678] <= 32'b001111_11110_01001_1111111111111101; 	// lw
disk[679] <= 32'b000000_01000_01001_01111_00000_000010; 	// mul
disk[680] <= 32'b001110_01111_00001_0000000000000000; 	// mov
disk[681] <= 32'b011010_00000_00001_0000000000000000; 	// mmuLowerIM
disk[682] <= 32'b010001_11101_01010_0000000011100011; 	// la
disk[683] <= 32'b001111_11110_01011_1111111111111001; 	// lw
disk[684] <= 32'b000000_01010_01011_10000_00000_000000; 	// add
disk[685] <= 32'b010010_10000_00111_0000000000000000; 	// sw
disk[686] <= 32'b010001_11101_01100_0000000011101101; 	// la
disk[687] <= 32'b000000_01100_01011_10001_00000_000000; 	// add
disk[688] <= 32'b001111_11110_01101_1111111111111111; 	// lw
disk[689] <= 32'b010010_10001_01101_0000000000000000; 	// sw
disk[690] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[691] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[692] <= 32'b010010_11110_00001_0000000000000000; 	// sw
disk[693] <= 32'b010001_11101_00101_0000000011100011; 	// la
disk[694] <= 32'b001111_11101_00110_0000000001000001; 	// lw
disk[695] <= 32'b000000_00101_00110_01111_00000_000000; 	// add
disk[696] <= 32'b001111_01111_01111_0000000000000000; 	// lw
disk[697] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[698] <= 32'b000000_01111_10001_10000_00000_001101; 	// ne
disk[699] <= 32'b010101_10000_00000_0000001011011110; 	// jf
disk[700] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[701] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[702] <= 32'b100100_00000_00001_0000000000000000; 	// lcdCurr
disk[703] <= 32'b001111_11101_01000_0000000100000001; 	// lw
disk[704] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[705] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[706] <= 32'b001110_11110_10010_0000000000000000; 	// mov
disk[707] <= 32'b000001_10010_10011_0000000000000001; 	// addi
disk[708] <= 32'b010010_11101_10011_0000000010001000; 	// sw
disk[709] <= 32'b010001_11101_01001_0000000000000100; 	// la
disk[710] <= 32'b000000_01001_00110_10100_00000_000000; 	// add
disk[711] <= 32'b001111_11101_01010_0000000000000000; 	// lw
disk[712] <= 32'b010010_10100_01010_0000000000000000; 	// sw
disk[713] <= 32'b010001_11101_01011_0000000000001110; 	// la
disk[714] <= 32'b000000_01011_00110_10101_00000_000000; 	// add
disk[715] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[716] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[717] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[718] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
disk[719] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[720] <= 32'b100000_00000000000000000000000000; 	// exec
disk[721] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[722] <= 32'b010001_11101_00101_0000000000000100; 	// la
disk[723] <= 32'b001111_11101_00110_0000000001000001; 	// lw
disk[724] <= 32'b000000_00101_00110_10111_00000_000000; 	// add
disk[725] <= 32'b010000_00000_11000_0000000000000000; 	// li
disk[726] <= 32'b010010_10111_11000_0000000000000000; 	// sw
disk[727] <= 32'b010001_11101_00111_0000000000001110; 	// la
disk[728] <= 32'b000000_00111_00110_01111_00000_000000; 	// add
disk[729] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[730] <= 32'b010010_01111_10000_0000000000000000; 	// sw
disk[731] <= 32'b001111_11101_01000_0000000011111010; 	// lw
disk[732] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[733] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[734] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[735] <= 32'b000001_11110_11110_0000000000001000; 	// addi
disk[736] <= 32'b010010_11110_00001_1111111111111011; 	// sw
disk[737] <= 32'b001111_11110_00101_1111111111111011; 	// lw
disk[738] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[739] <= 32'b100100_00000_00001_0000000000000000; 	// lcdCurr
disk[740] <= 32'b001111_11101_00110_0000000100000001; 	// lw
disk[741] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[742] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[743] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[744] <= 32'b001111_11101_01000_0000000001000001; 	// lw
disk[745] <= 32'b000000_00111_01000_01111_00000_000000; 	// add
disk[746] <= 32'b001111_11101_01001_0000000000000000; 	// lw
disk[747] <= 32'b010010_01111_01001_0000000000000000; 	// sw
disk[748] <= 32'b010001_11101_01010_0000000000110110; 	// la
disk[749] <= 32'b000000_01010_01000_10000_00000_000000; 	// add
disk[750] <= 32'b001111_10000_10000_0000000000000000; 	// lw
disk[751] <= 32'b010010_11110_10000_1111111111111101; 	// sw
disk[752] <= 32'b001110_11110_10001_0000000000000000; 	// mov
disk[753] <= 32'b000001_10001_10010_0000000000000001; 	// addi
disk[754] <= 32'b010010_11110_10010_1111111111111110; 	// sw
disk[755] <= 32'b001111_11110_01011_1111111111111101; 	// lw
disk[756] <= 32'b001111_11101_01100_0000000010000010; 	// lw
disk[757] <= 32'b000000_01011_01100_10011_00000_000010; 	// mul
disk[758] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[759] <= 32'b010001_11101_01101_0000000000101100; 	// la
disk[760] <= 32'b000000_01101_01000_10100_00000_000000; 	// add
disk[761] <= 32'b001111_10100_10100_0000000000000000; 	// lw
disk[762] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[763] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[764] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[765] <= 32'b000000_00101_10110_10101_00000_010000; 	// gt
disk[766] <= 32'b010101_10101_00000_0000001100010010; 	// jf
disk[767] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[768] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[769] <= 32'b001111_00001_10111_0000000000000000; 	// lw
disk[770] <= 32'b010010_11110_10111_1111111111111100; 	// sw
disk[771] <= 32'b001111_11110_00111_1111111111111100; 	// lw
disk[772] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[773] <= 32'b001111_11110_01000_1111111111111110; 	// lw
disk[774] <= 32'b001110_01000_00010_0000000000000000; 	// mov
disk[775] <= 32'b010010_00010_00001_0000000000000000; 	// sw
disk[776] <= 32'b000001_01000_11000_0000000000000001; 	// addi
disk[777] <= 32'b010010_11110_11000_1111111111111110; 	// sw
disk[778] <= 32'b001111_11110_01000_1111111111111110; 	// lw
disk[779] <= 32'b000001_00110_01111_0000000000000001; 	// addi
disk[780] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[781] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[782] <= 32'b000010_00101_10000_0000000000000001; 	// subi
disk[783] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[784] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[785] <= 32'b111100_00000000000000001011111011; 	// j
disk[786] <= 32'b001110_11110_10001_0000000000000000; 	// mov
disk[787] <= 32'b010001_11101_00101_0000000000101100; 	// la
disk[788] <= 32'b001111_11101_00110_0000000001000001; 	// lw
disk[789] <= 32'b000000_00101_00110_10010_00000_000000; 	// add
disk[790] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[791] <= 32'b000000_10001_10010_10011_00000_000000; 	// add
disk[792] <= 32'b001110_10011_00001_0000000000000000; 	// mov
disk[793] <= 32'b001110_00001_11100_0000000000000000; 	// mov
disk[794] <= 32'b000001_00110_10100_0000000000000001; 	// addi
disk[795] <= 32'b001110_10100_00001_0000000000000000; 	// mov
disk[796] <= 32'b010001_11101_00111_0000000000001110; 	// la
disk[797] <= 32'b000000_00111_00110_10101_00000_000000; 	// add
disk[798] <= 32'b001111_10101_10101_0000000000000000; 	// lw
disk[799] <= 32'b001110_10101_00010_0000000000000000; 	// mov
disk[800] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
disk[801] <= 32'b010010_11110_11111_1111111111111010; 	// sw
disk[802] <= 32'b001110_11100_11110_0000000000000000; 	// mov
disk[803] <= 32'b001110_11011_11101_0000000000000000; 	// mov
disk[804] <= 32'b001110_00010_11010_0000000000000000; 	// mov
disk[805] <= 32'b001111_00000_00000_0000011111100000; 	// lw
disk[806] <= 32'b001111_00000_00001_0000011111100001; 	// lw
disk[807] <= 32'b001111_00000_00010_0000011111100010; 	// lw
disk[808] <= 32'b001111_00000_00011_0000011111100011; 	// lw
disk[809] <= 32'b001111_00000_00100_0000011111100100; 	// lw
disk[810] <= 32'b001111_00000_00101_0000011111100101; 	// lw
disk[811] <= 32'b001111_00000_00110_0000011111100110; 	// lw
disk[812] <= 32'b001111_00000_00111_0000011111100111; 	// lw
disk[813] <= 32'b001111_00000_01000_0000011111101000; 	// lw
disk[814] <= 32'b001111_00000_01001_0000011111101001; 	// lw
disk[815] <= 32'b001111_00000_01010_0000011111101010; 	// lw
disk[816] <= 32'b001111_00000_01011_0000011111101011; 	// lw
disk[817] <= 32'b001111_00000_01100_0000011111101100; 	// lw
disk[818] <= 32'b001111_00000_01101_0000011111101101; 	// lw
disk[819] <= 32'b001111_00000_01110_0000011111101110; 	// lw
disk[820] <= 32'b001111_00000_01111_0000011111101111; 	// lw
disk[821] <= 32'b001111_00000_10000_0000011111110000; 	// lw
disk[822] <= 32'b001111_00000_10001_0000011111110001; 	// lw
disk[823] <= 32'b001111_00000_10010_0000011111110010; 	// lw
disk[824] <= 32'b001111_00000_10011_0000011111110011; 	// lw
disk[825] <= 32'b001111_00000_10100_0000011111110100; 	// lw
disk[826] <= 32'b001111_00000_10101_0000011111110101; 	// lw
disk[827] <= 32'b001111_00000_10110_0000011111110110; 	// lw
disk[828] <= 32'b001111_00000_10111_0000011111110111; 	// lw
disk[829] <= 32'b001111_00000_11000_0000011111111000; 	// lw
disk[830] <= 32'b001111_00000_11001_0000011111111001; 	// lw
disk[831] <= 32'b100001_11010_00000_0000000000000000; 	// execAgain
disk[832] <= 32'b001111_11110_11111_1111111111111010; 	// lw
disk[833] <= 32'b010001_11101_00101_0000000000000100; 	// la
disk[834] <= 32'b001111_11101_00110_0000000001000001; 	// lw
disk[835] <= 32'b000000_00101_00110_10110_00000_000000; 	// add
disk[836] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[837] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[838] <= 32'b010001_11101_00111_0000000000001110; 	// la
disk[839] <= 32'b000000_00111_00110_11000_00000_000000; 	// add
disk[840] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[841] <= 32'b010010_11000_01111_0000000000000000; 	// sw
disk[842] <= 32'b001111_11101_01000_0000000011111010; 	// lw
disk[843] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[844] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[845] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[846] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[847] <= 32'b010010_11110_00001_0000000000000000; 	// sw
disk[848] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[849] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[850] <= 32'b010010_11101_01111_0000000001000001; 	// sw
disk[851] <= 32'b001111_11101_00110_0000000001000001; 	// lw
disk[852] <= 32'b010010_11101_00110_0000000001000000; 	// sw
disk[853] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[854] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[855] <= 32'b111110_00000000000000001010110011; 	// jal
disk[856] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[857] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[858] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[859] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[860] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[861] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[862] <= 32'b111110_00000000000000001000101111; 	// jal
disk[863] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[864] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[865] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[866] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[867] <= 32'b111110_00000000000000001000011000; 	// jal
disk[868] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[869] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[870] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[871] <= 32'b001111_11101_00110_0000000000000011; 	// lw
disk[872] <= 32'b000000_00101_00110_01111_00000_001101; 	// ne
disk[873] <= 32'b010101_01111_00000_0000001101111001; 	// jf
disk[874] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[875] <= 32'b111110_00000000000000001000011000; 	// jal
disk[876] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[877] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[878] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[879] <= 32'b010010_11101_00101_0000000001000001; 	// sw
disk[880] <= 32'b001111_11101_00110_0000000001000001; 	// lw
disk[881] <= 32'b000001_00110_10000_0000000000000001; 	// addi
disk[882] <= 32'b001110_10000_00001_0000000000000000; 	// mov
disk[883] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[884] <= 32'b111110_00000000000000001010110011; 	// jal
disk[885] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[886] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[887] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[888] <= 32'b111100_00000000000000001101100010; 	// j
disk[889] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[890] <= 32'b001110_11110_11100_0000000000000000; 	// mov
disk[891] <= 32'b001110_11101_11011_0000000000000000; 	// mov
disk[892] <= 32'b010000_00000_00000_0000000000000000; 	// li
disk[893] <= 32'b010000_00000_11110_0000000000000000; 	// li
disk[894] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[895] <= 32'b000001_11110_11110_0000000100001100; 	// addi
disk[896] <= 32'b010010_00000_00000_0000011111100000; 	// sw
disk[897] <= 32'b010010_00000_00001_0000011111100001; 	// sw
disk[898] <= 32'b010010_00000_00010_0000011111100010; 	// sw
disk[899] <= 32'b010010_00000_00011_0000011111100011; 	// sw
disk[900] <= 32'b010010_00000_00100_0000011111100100; 	// sw
disk[901] <= 32'b010010_00000_00101_0000011111100101; 	// sw
disk[902] <= 32'b010010_00000_00110_0000011111100110; 	// sw
disk[903] <= 32'b010010_00000_00111_0000011111100111; 	// sw
disk[904] <= 32'b010010_00000_01000_0000011111101000; 	// sw
disk[905] <= 32'b010010_00000_01001_0000011111101001; 	// sw
disk[906] <= 32'b010010_00000_01010_0000011111101010; 	// sw
disk[907] <= 32'b010010_00000_01011_0000011111101011; 	// sw
disk[908] <= 32'b010010_00000_01100_0000011111101100; 	// sw
disk[909] <= 32'b010010_00000_01101_0000011111101101; 	// sw
disk[910] <= 32'b010010_00000_01110_0000011111101110; 	// sw
disk[911] <= 32'b010010_00000_01111_0000011111101111; 	// sw
disk[912] <= 32'b010010_00000_10000_0000011111110000; 	// sw
disk[913] <= 32'b010010_00000_10001_0000011111110001; 	// sw
disk[914] <= 32'b010010_00000_10010_0000011111110010; 	// sw
disk[915] <= 32'b010010_00000_10011_0000011111110011; 	// sw
disk[916] <= 32'b010010_00000_10100_0000011111110100; 	// sw
disk[917] <= 32'b010010_00000_10101_0000011111110101; 	// sw
disk[918] <= 32'b010010_00000_10110_0000011111110110; 	// sw
disk[919] <= 32'b010010_00000_10111_0000011111110111; 	// sw
disk[920] <= 32'b010010_00000_11000_0000011111111000; 	// sw
disk[921] <= 32'b010010_00000_11001_0000011111111001; 	// sw
disk[922] <= 32'b001111_11110_00101_1111111111111011; 	// lw
disk[923] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[924] <= 32'b000000_00101_10000_01111_00000_001100; 	// eq
disk[925] <= 32'b010101_01111_00000_0000001110100111; 	// jf
disk[926] <= 32'b111110_00000000000000000100101101; 	// jal
disk[927] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[928] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[929] <= 32'b001111_11101_00110_0000000011111010; 	// lw
disk[930] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[931] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[932] <= 32'b010000_00000_10001_0000000000000001; 	// li
disk[933] <= 32'b010010_11110_10001_1111111111111011; 	// sw
disk[934] <= 32'b100110_00000_00000_0000000000000000; 	// cic
disk[935] <= 32'b100101_00000_10010_0000000000000000; 	// gic
disk[936] <= 32'b010010_11110_10010_1111111111111010; 	// sw
disk[937] <= 32'b001111_11110_00101_1111111111111010; 	// lw
disk[938] <= 32'b010000_00000_10100_0000000000000001; 	// li
disk[939] <= 32'b000000_00101_10100_10011_00000_001100; 	// eq
disk[940] <= 32'b010101_10011_00000_0000010000100111; 	// jf
disk[941] <= 32'b001110_11100_10101_0000000000000000; 	// mov
disk[942] <= 32'b010010_11101_10101_0000000010001001; 	// sw
disk[943] <= 32'b001111_11101_00110_0000000010001001; 	// lw
disk[944] <= 32'b001111_11101_00111_0000000010001000; 	// lw
disk[945] <= 32'b000000_00110_00111_10110_00000_000001; 	// sub
disk[946] <= 32'b000001_10110_10111_0000000000000001; 	// addi
disk[947] <= 32'b010010_11110_10111_0000000000000000; 	// sw
disk[948] <= 32'b010001_11101_01000_0000000000101100; 	// la
disk[949] <= 32'b001111_11101_01001_0000000001000001; 	// lw
disk[950] <= 32'b000000_01000_01001_11000_00000_000000; 	// add
disk[951] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[952] <= 32'b010010_11000_01010_0000000000000000; 	// sw
disk[953] <= 32'b010001_11101_01011_0000000000000100; 	// la
disk[954] <= 32'b000000_01011_01001_01111_00000_000000; 	// add
disk[955] <= 32'b001111_11101_01100_0000000000000010; 	// lw
disk[956] <= 32'b010010_01111_01100_0000000000000000; 	// sw
disk[957] <= 32'b100111_00000_10000_0000000000000000; 	// gip
disk[958] <= 32'b000001_10000_10001_0000000000000001; 	// addi
disk[959] <= 32'b010001_11101_01101_0000000000001110; 	// la
disk[960] <= 32'b000000_01101_01001_10010_00000_000000; 	// add
disk[961] <= 32'b010010_10010_10001_0000000000000000; 	// sw
disk[962] <= 32'b010001_11101_01110_0000000000110110; 	// la
disk[963] <= 32'b000000_01110_01001_10011_00000_000000; 	// add
disk[964] <= 32'b001111_10011_10011_0000000000000000; 	// lw
disk[965] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[966] <= 32'b000000_10011_10101_10100_00000_001100; 	// eq
disk[967] <= 32'b010101_10100_00000_0000001111010010; 	// jf
disk[968] <= 32'b111110_00000000000000000110000011; 	// jal
disk[969] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[970] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[971] <= 32'b010010_11110_00101_1111111111111100; 	// sw
disk[972] <= 32'b010001_11101_00110_0000000000110110; 	// la
disk[973] <= 32'b001111_11101_00111_0000000001000001; 	// lw
disk[974] <= 32'b000000_00110_00111_10110_00000_000000; 	// add
disk[975] <= 32'b001111_11110_01000_1111111111111100; 	// lw
disk[976] <= 32'b010010_10110_01000_0000000000000000; 	// sw
disk[977] <= 32'b111100_00000000000000001111010111; 	// j
disk[978] <= 32'b010001_11101_00101_0000000000110110; 	// la
disk[979] <= 32'b001111_11101_00110_0000000001000001; 	// lw
disk[980] <= 32'b000000_00101_00110_10111_00000_000000; 	// add
disk[981] <= 32'b001111_10111_10111_0000000000000000; 	// lw
disk[982] <= 32'b010010_11110_10111_1111111111111100; 	// sw
disk[983] <= 32'b001111_11101_00101_0000000010001000; 	// lw
disk[984] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[985] <= 32'b001111_11110_00110_1111111111111100; 	// lw
disk[986] <= 32'b001111_11101_00111_0000000010000010; 	// lw
disk[987] <= 32'b000000_00110_00111_11000_00000_000010; 	// mul
disk[988] <= 32'b010010_11110_11000_1111111111111111; 	// sw
disk[989] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[990] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[991] <= 32'b000000_00101_10000_01111_00000_010000; 	// gt
disk[992] <= 32'b010101_01111_00000_0000001111110100; 	// jf
disk[993] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[994] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[995] <= 32'b001111_00001_10001_0000000000000000; 	// lw
disk[996] <= 32'b010010_11110_10001_1111111111111101; 	// sw
disk[997] <= 32'b001111_11110_00111_1111111111111101; 	// lw
disk[998] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[999] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[1000] <= 32'b001110_01000_00010_0000000000000000; 	// mov
disk[1001] <= 32'b010010_00010_00001_0000000000000000; 	// sw
disk[1002] <= 32'b000001_00110_10010_0000000000000001; 	// addi
disk[1003] <= 32'b010010_11110_10010_1111111111111110; 	// sw
disk[1004] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[1005] <= 32'b000001_01000_10011_0000000000000001; 	// addi
disk[1006] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[1007] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[1008] <= 32'b000010_00101_10100_0000000000000001; 	// subi
disk[1009] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[1010] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1011] <= 32'b111100_00000000000000001111011101; 	// j
disk[1012] <= 32'b001111_11101_00101_0000000001000001; 	// lw
disk[1013] <= 32'b001111_11101_00110_0000000001000000; 	// lw
disk[1014] <= 32'b000000_00101_00110_10101_00000_001100; 	// eq
disk[1015] <= 32'b010101_10101_00000_0000010000000001; 	// jf
disk[1016] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1017] <= 32'b111110_00000000000000001011011111; 	// jal
disk[1018] <= 32'b000010_11110_11110_0000000000001000; 	// subi
disk[1019] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[1020] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[1021] <= 32'b010000_00000_11110_0000000100001100; 	// li
disk[1022] <= 32'b010000_00000_10110_0000001111100111; 	// li
disk[1023] <= 32'b010010_11101_10110_0000000001000000; 	// sw
disk[1024] <= 32'b111100_00000000000000010000100001; 	// j
disk[1025] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[1026] <= 32'b000001_00101_10111_0000000000000001; 	// addi
disk[1027] <= 32'b010010_11110_10111_1111111111111100; 	// sw
disk[1028] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[1029] <= 32'b001111_11101_00110_0000000010000011; 	// lw
disk[1030] <= 32'b000010_00110_11000_0000000000000001; 	// subi
disk[1031] <= 32'b001111_11101_00111_0000000010000010; 	// lw
disk[1032] <= 32'b000000_00111_11000_01111_00000_000010; 	// mul
disk[1033] <= 32'b010010_11110_01111_1111111111111110; 	// sw
disk[1034] <= 32'b000000_00101_00111_10000_00000_000010; 	// mul
disk[1035] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[1036] <= 32'b001111_11101_00101_0000000010000010; 	// lw
disk[1037] <= 32'b001111_11101_00110_0000000010000011; 	// lw
disk[1038] <= 32'b000000_00101_00110_10001_00000_000010; 	// mul
disk[1039] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[1040] <= 32'b000000_00111_10001_10010_00000_001110; 	// lt
disk[1041] <= 32'b010101_10010_00000_0000010000100001; 	// jf
disk[1042] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1043] <= 32'b001111_00001_10011_0000000000000000; 	// lw
disk[1044] <= 32'b010010_11110_10011_1111111111111101; 	// sw
disk[1045] <= 32'b001111_11110_01000_1111111111111101; 	// lw
disk[1046] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[1047] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[1048] <= 32'b001110_01001_00010_0000000000000000; 	// mov
disk[1049] <= 32'b010010_00010_00001_0000000000000000; 	// sw
disk[1050] <= 32'b000001_00111_10100_0000000000000001; 	// addi
disk[1051] <= 32'b010010_11110_10100_1111111111111110; 	// sw
disk[1052] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[1053] <= 32'b000001_01001_10101_0000000000000001; 	// addi
disk[1054] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[1055] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[1056] <= 32'b111100_00000000000000010000001100; 	// j
disk[1057] <= 32'b001111_11101_00101_0000000011111010; 	// lw
disk[1058] <= 32'b010010_11101_00101_0000000100000010; 	// sw
disk[1059] <= 32'b001111_11101_00110_0000000100000010; 	// lw
disk[1060] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1061] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[1062] <= 32'b100110_00000_00000_0000000000000000; 	// cic
disk[1063] <= 32'b010000_00000_10110_0000000000000001; 	// li
disk[1064] <= 32'b010101_10110_00000_0000010011001100; 	// jf
disk[1065] <= 32'b010011_00000_10111_0000000000000000; 	// in
disk[1066] <= 32'b010010_11110_10111_1111111111111001; 	// sw
disk[1067] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1068] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1069] <= 32'b010000_00000_00010_0000000000000000; 	// li
disk[1070] <= 32'b010100_00000_00001_0000000000000000; 	// out
disk[1071] <= 32'b001111_11101_00110_0000000100000010; 	// lw
disk[1072] <= 32'b001111_11101_00111_0000000011111010; 	// lw
disk[1073] <= 32'b000000_00110_00111_11000_00000_001100; 	// eq
disk[1074] <= 32'b010101_11000_00000_0000010001001011; 	// jf
disk[1075] <= 32'b010000_00000_10000_0000000000000100; 	// li
disk[1076] <= 32'b000000_00101_10000_01111_00000_010000; 	// gt
disk[1077] <= 32'b010101_01111_00000_0000010000111001; 	// jf
disk[1078] <= 32'b010010_11110_00111_1111111111111001; 	// sw
disk[1079] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1080] <= 32'b111100_00000000000000010001001010; 	// j
disk[1081] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1082] <= 32'b010000_00000_10010_0000000000000100; 	// li
disk[1083] <= 32'b000000_00101_10010_10001_00000_001100; 	// eq
disk[1084] <= 32'b010101_10001_00000_0000010001000011; 	// jf
disk[1085] <= 32'b111110_00000000000000000000110011; 	// jal
disk[1086] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[1087] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[1088] <= 32'b001111_11101_00110_0000000011111010; 	// lw
disk[1089] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1090] <= 32'b111100_00000000000000010001001010; 	// j
disk[1091] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1092] <= 32'b010000_00000_10100_0000000000000001; 	// li
disk[1093] <= 32'b000000_00101_10100_10011_00000_001110; 	// lt
disk[1094] <= 32'b010101_10011_00000_0000010001001010; 	// jf
disk[1095] <= 32'b001111_11101_00110_0000000011111010; 	// lw
disk[1096] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1097] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1098] <= 32'b111100_00000000000000010011000110; 	// j
disk[1099] <= 32'b001111_11101_00101_0000000100000010; 	// lw
disk[1100] <= 32'b001111_11101_00110_0000000011111011; 	// lw
disk[1101] <= 32'b000000_00101_00110_10101_00000_001100; 	// eq
disk[1102] <= 32'b010101_10101_00000_0000010001011111; 	// jf
disk[1103] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1104] <= 32'b010000_00000_10111_0000000000000011; 	// li
disk[1105] <= 32'b000000_00111_10111_10110_00000_010000; 	// gt
disk[1106] <= 32'b010101_10110_00000_0000010001010111; 	// jf
disk[1107] <= 32'b001111_11101_01000_0000000011111010; 	// lw
disk[1108] <= 32'b010010_11110_01000_1111111111111001; 	// sw
disk[1109] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1110] <= 32'b111100_00000000000000010001011110; 	// j
disk[1111] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1112] <= 32'b010000_00000_01111_0000000000000001; 	// li
disk[1113] <= 32'b000000_00101_01111_11000_00000_001110; 	// lt
disk[1114] <= 32'b010101_11000_00000_0000010001011110; 	// jf
disk[1115] <= 32'b001111_11101_00110_0000000011111010; 	// lw
disk[1116] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1117] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1118] <= 32'b111100_00000000000000010011000110; 	// j
disk[1119] <= 32'b001111_11101_00101_0000000100000010; 	// lw
disk[1120] <= 32'b001111_11101_00110_0000000011111100; 	// lw
disk[1121] <= 32'b000000_00101_00110_10000_00000_001100; 	// eq
disk[1122] <= 32'b010101_10000_00000_0000010010000000; 	// jf
disk[1123] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1124] <= 32'b010000_00000_10010_0000000000000001; 	// li
disk[1125] <= 32'b000000_00111_10010_10001_00000_001100; 	// eq
disk[1126] <= 32'b010101_10001_00000_0000010001110000; 	// jf
disk[1127] <= 32'b001111_11101_01000_0000000011111110; 	// lw
disk[1128] <= 32'b010010_11110_01000_1111111111111001; 	// sw
disk[1129] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1130] <= 32'b111110_00000000000000000111100000; 	// jal
disk[1131] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1132] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[1133] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1134] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[1135] <= 32'b111100_00000000000000010001111111; 	// j
disk[1136] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1137] <= 32'b010000_00000_10100_0000000000000011; 	// li
disk[1138] <= 32'b000000_00101_10100_10011_00000_010000; 	// gt
disk[1139] <= 32'b010101_10011_00000_0000010001111000; 	// jf
disk[1140] <= 32'b001111_11101_00110_0000000011111010; 	// lw
disk[1141] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1142] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1143] <= 32'b111100_00000000000000010001111111; 	// j
disk[1144] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1145] <= 32'b010000_00000_10110_0000000000000001; 	// li
disk[1146] <= 32'b000000_00101_10110_10101_00000_001110; 	// lt
disk[1147] <= 32'b010101_10101_00000_0000010001111111; 	// jf
disk[1148] <= 32'b001111_11101_00110_0000000011111010; 	// lw
disk[1149] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1150] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1151] <= 32'b111100_00000000000000010011000110; 	// j
disk[1152] <= 32'b001111_11101_00101_0000000100000010; 	// lw
disk[1153] <= 32'b001111_11101_00110_0000000011111101; 	// lw
disk[1154] <= 32'b000000_00101_00110_10111_00000_001100; 	// eq
disk[1155] <= 32'b010101_10111_00000_0000010010101001; 	// jf
disk[1156] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1157] <= 32'b010000_00000_01111_0000000000000001; 	// li
disk[1158] <= 32'b000000_00111_01111_11000_00000_001100; 	// eq
disk[1159] <= 32'b010101_11000_00000_0000010010001110; 	// jf
disk[1160] <= 32'b111110_00000000000000001101011100; 	// jal
disk[1161] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[1162] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[1163] <= 32'b001111_11101_00110_0000000011111010; 	// lw
disk[1164] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1165] <= 32'b111100_00000000000000010010101000; 	// j
disk[1166] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1167] <= 32'b010000_00000_10001_0000000000000010; 	// li
disk[1168] <= 32'b000000_00101_10001_10000_00000_001100; 	// eq
disk[1169] <= 32'b010101_10000_00000_0000010010011010; 	// jf
disk[1170] <= 32'b111110_00000000000000000110111111; 	// jal
disk[1171] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1172] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[1173] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1174] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[1175] <= 32'b001111_11101_00110_0000000011111111; 	// lw
disk[1176] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1177] <= 32'b111100_00000000000000010010101000; 	// j
disk[1178] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1179] <= 32'b010000_00000_10011_0000000000000011; 	// li
disk[1180] <= 32'b000000_00101_10011_10010_00000_001100; 	// eq
disk[1181] <= 32'b010101_10010_00000_0000010010100110; 	// jf
disk[1182] <= 32'b111110_00000000000000000110111111; 	// jal
disk[1183] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1184] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[1185] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1186] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[1187] <= 32'b001111_11101_00110_0000000100000000; 	// lw
disk[1188] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1189] <= 32'b111100_00000000000000010010101000; 	// j
disk[1190] <= 32'b001111_11101_00101_0000000011111010; 	// lw
disk[1191] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1192] <= 32'b111100_00000000000000010011000110; 	// j
disk[1193] <= 32'b001111_11101_00101_0000000100000010; 	// lw
disk[1194] <= 32'b001111_11101_00110_0000000011111110; 	// lw
disk[1195] <= 32'b000000_00101_00110_10100_00000_001100; 	// eq
disk[1196] <= 32'b010101_10100_00000_0000010010111000; 	// jf
disk[1197] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1198] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[1199] <= 32'b000000_00111_10110_10101_00000_010000; 	// gt
disk[1200] <= 32'b010101_10101_00000_0000010010110101; 	// jf
disk[1201] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1202] <= 32'b111110_00000000000000001001100001; 	// jal
disk[1203] <= 32'b000010_11110_11110_0000000000001010; 	// subi
disk[1204] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[1205] <= 32'b001111_11101_00101_0000000011111010; 	// lw
disk[1206] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1207] <= 32'b111100_00000000000000010011000110; 	// j
disk[1208] <= 32'b001111_11101_00101_0000000100000010; 	// lw
disk[1209] <= 32'b001111_11101_00110_0000000011111111; 	// lw
disk[1210] <= 32'b000000_00101_00110_10111_00000_001100; 	// eq
disk[1211] <= 32'b010101_10111_00000_0000010011000110; 	// jf
disk[1212] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1213] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[1214] <= 32'b000000_00111_01111_11000_00000_010000; 	// gt
disk[1215] <= 32'b010101_11000_00000_0000010011000100; 	// jf
disk[1216] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1217] <= 32'b111110_00000000000000001101001110; 	// jal
disk[1218] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1219] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[1220] <= 32'b001111_11101_00101_0000000011111010; 	// lw
disk[1221] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1222] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1223] <= 32'b010010_11101_00101_0000000100000010; 	// sw
disk[1224] <= 32'b001111_11101_00110_0000000100000010; 	// lw
disk[1225] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1226] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[1227] <= 32'b111100_00000000000000010000100111; 	// j
disk[1228] <= 32'b111111_00000000000000000000000000; 	// halt

		// PROGRAMA 1
		disk[1700] <= 32'b111101_00000000000000000000100011;		// Jump to Main
		disk[1701] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[1702] <= 32'b010010_11110_00001_1111111111111100; 	// sw
		disk[1703] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[1704] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[1705] <= 32'b010000_00000_10000_0000000000000001; 	// li
		disk[1706] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[1707] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[1708] <= 32'b010010_11110_10001_1111111111111101; 	// sw
		disk[1709] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[1710] <= 32'b001111_11110_00110_1111111111111100; 	// lw
		disk[1711] <= 32'b000000_00101_00110_10010_00000_001111; 	// let
		disk[1712] <= 32'b010101_10010_00000_0000000000100000; 	// jf
		disk[1713] <= 32'b010000_00000_10100_0000000000000001; 	// li
		disk[1714] <= 32'b000000_00101_10100_10011_00000_001111; 	// let
		disk[1715] <= 32'b010101_10011_00000_0000000000010010; 	// jf
		disk[1716] <= 32'b010010_11110_00101_1111111111111110; 	// sw
		disk[1717] <= 32'b111100_00000000000000000000011011; 	// j
		disk[1718] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1719] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[1720] <= 32'b000000_00101_00110_10101_00000_000000; 	// add
		disk[1721] <= 32'b010010_11110_10101_1111111111111110; 	// sw
		disk[1722] <= 32'b010010_11110_00110_1111111111111111; 	// sw
		disk[1723] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1724] <= 32'b001111_11110_00111_1111111111111110; 	// lw
		disk[1725] <= 32'b010010_11110_00111_0000000000000000; 	// sw
		disk[1726] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[1727] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[1728] <= 32'b000001_00101_10110_0000000000000001; 	// addi
		disk[1729] <= 32'b010010_11110_10110_1111111111111101; 	// sw
		disk[1730] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[1731] <= 32'b111100_00000000000000000000001001; 	// j
		disk[1732] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[1733] <= 32'b001110_00101_11001_0000000000000000; 	// mov
		disk[1734] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1735] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[1736] <= 32'b010000_00000_01111_0000000000001011; 	// li
		disk[1737] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[1738] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1739] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1740] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1741] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[1742] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[1743] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1744] <= 32'b001110_11001_00101_0000000000000000; 	// mov
		disk[1745] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1746] <= 32'b010000_00000_00010_0000000000000000; 	// li
		disk[1747] <= 32'b010100_00000_00001_0000000000000000; 	// out
		disk[1748] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[1749] <= 32'b011111_11111_00000_0000000000000000; 	// syscall

		// PROGRAMA 2
		disk[1800] <= 32'b111101_00000000000000000000100001;		// Jump to Main
		disk[1801] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[1802] <= 32'b010010_11110_00001_1111111111111100; 	// sw
		disk[1803] <= 32'b010010_11110_00010_1111111111111101; 	// sw
		disk[1804] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[1805] <= 32'b010010_11110_01111_1111111111111110; 	// sw
		disk[1806] <= 32'b010000_00000_10000_0000000000000000; 	// li
		disk[1807] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[1808] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[1809] <= 32'b001111_11110_00110_1111111111111101; 	// lw
		disk[1810] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
		disk[1811] <= 32'b010101_10001_00000_0000000000011100; 	// jf
		disk[1812] <= 32'b001111_11110_00111_1111111111111100; 	// lw
		disk[1813] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
		disk[1814] <= 32'b001111_10010_10010_0000000000000000; 	// lw
		disk[1815] <= 32'b001111_11110_01000_0000000000000000; 	// lw
		disk[1816] <= 32'b000000_01000_10010_10011_00000_001110; 	// lt
		disk[1817] <= 32'b010101_10011_00000_0000000000010111; 	// jf
		disk[1818] <= 32'b000000_00111_00101_10100_00000_000000; 	// add
		disk[1819] <= 32'b001111_10100_10100_0000000000000000; 	// lw
		disk[1820] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[1821] <= 32'b001111_11110_01000_0000000000000000; 	// lw
		disk[1822] <= 32'b010010_11110_00101_1111111111111111; 	// sw
		disk[1823] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[1824] <= 32'b000001_00101_10101_0000000000000001; 	// addi
		disk[1825] <= 32'b010010_11110_10101_1111111111111110; 	// sw
		disk[1826] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[1827] <= 32'b111100_00000000000000000000001000; 	// j
		disk[1828] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1829] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1830] <= 32'b010000_00000_00010_0000000000000001; 	// li
		disk[1831] <= 32'b010100_00000_00001_0000000000000001; 	// out
		disk[1832] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1833] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[1834] <= 32'b010001_11110_00101_1111111111111011; 	// la
		disk[1835] <= 32'b010000_00000_01111_0000000000001100; 	// li
		disk[1836] <= 32'b010010_00101_01111_0000000000000000; 	// sw
		disk[1837] <= 32'b010000_00000_10000_0000000000101001; 	// li
		disk[1838] <= 32'b010010_00101_10000_0000000000000001; 	// sw
		disk[1839] <= 32'b010000_00000_10001_0000000000010111; 	// li
		disk[1840] <= 32'b010010_00101_10001_0000000000000010; 	// sw
		disk[1841] <= 32'b010000_00000_10010_0000000001100010; 	// li
		disk[1842] <= 32'b010010_00101_10010_0000000000000011; 	// sw
		disk[1843] <= 32'b010000_00000_10011_0000000000100001; 	// li
		disk[1844] <= 32'b010010_00101_10011_0000000000000100; 	// sw
		disk[1845] <= 32'b010000_00000_10100_0000000000010101; 	// li
		disk[1846] <= 32'b010010_00101_10100_0000000000000101; 	// sw
		disk[1847] <= 32'b010001_11110_00001_1111111111111011; 	// la
		disk[1848] <= 32'b010000_00000_00010_0000000000000110; 	// li
		disk[1849] <= 32'b010010_11110_11111_1111111111111010; 	// sw
		disk[1850] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[1851] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[1852] <= 32'b001111_11110_11111_1111111111111010; 	// lw
		disk[1853] <= 32'b001110_11001_00101_0000000000000000; 	// mov
		disk[1854] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[1855] <= 32'b011111_11111_00000_0000000000000000; 	// syscall
		
		// PROGRAMA 3
		disk[1900] <= 32'b111101_00000000000000000000010100;		// Jump to Main
		disk[1901] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[1902] <= 32'b010010_11110_00001_1111111111111111; 	// sw
		disk[1903] <= 32'b010000_00000_01111_0000000000000001; 	// li
		disk[1904] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[1905] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1906] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[1907] <= 32'b000000_00101_10001_10000_00000_010000; 	// gt
		disk[1908] <= 32'b010101_10000_00000_0000000000010001; 	// jf
		disk[1909] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[1910] <= 32'b000000_00110_00101_10010_00000_000010; 	// mul
		disk[1911] <= 32'b010010_11110_10010_0000000000000000; 	// sw
		disk[1912] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[1913] <= 32'b000010_00101_10011_0000000000000001; 	// subi
		disk[1914] <= 32'b010010_11110_10011_1111111111111111; 	// sw
		disk[1915] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1916] <= 32'b111100_00000000000000000000000101; 	// j
		disk[1917] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1918] <= 32'b001110_00101_11001_0000000000000000; 	// mov
		disk[1919] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1920] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[1921] <= 32'b010000_00000_01111_0000000001011101; 	// li
		disk[1922] <= 32'b010010_11110_01111_1111111111111110; 	// sw
		disk[1923] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[1924] <= 32'b010010_11110_00101_1111111111111111; 	// sw
		disk[1925] <= 32'b101000_00000000000000000000000000; 	// preIO
		disk[1926] <= 32'b010011_00000_10000_0000000000000000; 	// in
		disk[1927] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[1928] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1929] <= 32'b010000_00000_00010_0000000000000000; 	// li
		disk[1930] <= 32'b010100_00000_00001_0000000000000000; 	// out
		disk[1931] <= 32'b001111_11110_00110_1111111111111111; 	// lw
		disk[1932] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[1933] <= 32'b010000_00000_00010_0000000000000001; 	// li
		disk[1934] <= 32'b010100_00000_00001_0000000000000001; 	// out
		disk[1935] <= 32'b001111_11110_00111_0000000000000000; 	// lw
		disk[1936] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[1937] <= 32'b010010_11110_11111_1111111111111101; 	// sw
		disk[1938] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[1939] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[1940] <= 32'b001111_11110_11111_1111111111111101; 	// lw
		disk[1941] <= 32'b001110_11001_00101_0000000000000000; 	// mov
		disk[1942] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1943] <= 32'b010000_00000_00010_0000000000000010; 	// li
		disk[1944] <= 32'b010100_00000_00001_0000000000000010; 	// out
		disk[1945] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[1946] <= 32'b011111_11111_00000_0000000000000000; 	// syscall

	end
endmodule
