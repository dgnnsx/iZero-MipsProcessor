module disco_rigido (clk, we, addr, datain, dataout);
	input clk;										// clock
	input we;										// write enable
	input [31:0] addr;							// disk address
	input [31:0] datain;							// data in (to disk)
	
	output reg [31:0] dataout;					// data out (from disk)
	
	localparam DISK_SIZE = 2048;				// Tamanho do disco
	reg [31:0] disk [DISK_SIZE-1:0];			// disk cells
	
	always @ (posedge clk) begin
		if (we) disk[addr] <= datain;			// write disk
	end
	
	always @ (negedge clk) begin
		dataout <= disk[addr];
	end

	initial begin
		// SISTEMA OPERACIONAL

disk[0] <= 32'b111100_00000000000000001001010100;		// Jump to Main
disk[1] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[2] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[3] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[4] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[5] <= 32'b001110_01010_00110_0000000000000000; 	// mov
disk[6] <= 32'b010110_00110_10101_0000000000000000; 	// ldk
disk[7] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[8] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[9] <= 32'b001101_01010_10110_0000000000011010; 	// srli
disk[10] <= 32'b001111_00101_01011_0000000010011100; 	// lw
disk[11] <= 32'b000000_10110_01011_10111_00000_001101; 	// ne
disk[12] <= 32'b010101_10111_00000_0000000000010110; 	// jf
disk[13] <= 32'b001111_11110_01100_0000000000000000; 	// lw
disk[14] <= 32'b000001_01100_11000_0000000000000001; 	// addi
disk[15] <= 32'b010010_11110_11000_0000000000000000; 	// sw
disk[16] <= 32'b001111_11110_01100_0000000000000000; 	// lw
disk[17] <= 32'b001110_01100_00110_0000000000000000; 	// mov
disk[18] <= 32'b010110_00110_11001_0000000000000000; 	// ldk
disk[19] <= 32'b010010_11110_11001_1111111111111111; 	// sw
disk[20] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[21] <= 32'b111100_00000000000000000000001000; 	// j
disk[22] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[23] <= 32'b001110_01010_00001_0000000000000000; 	// mov
disk[24] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[25] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[26] <= 32'b010010_11110_00110_1111111111111111; 	// sw
disk[27] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[28] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[29] <= 32'b000000_01010_10101_10100_00000_001100; 	// eq
disk[30] <= 32'b010101_10100_00000_0000000000100010; 	// jf
disk[31] <= 32'b010000_00000_10110_0000000000000001; 	// li
disk[32] <= 32'b001110_10110_00001_0000000000000000; 	// mov
disk[33] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[34] <= 32'b010000_00000_10111_0000000000000001; 	// li
disk[35] <= 32'b010010_11110_10111_0000000000000000; 	// sw
disk[36] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[37] <= 32'b010000_00000_11001_0000000000000000; 	// li
disk[38] <= 32'b000000_01010_11001_11000_00000_010000; 	// gt
disk[39] <= 32'b010101_11000_00000_0000000000110000; 	// jf
disk[40] <= 32'b001111_11110_01011_0000000000000000; 	// lw
disk[41] <= 32'b000011_01011_11010_0000000000000010; 	// muli
disk[42] <= 32'b010010_11110_11010_0000000000000000; 	// sw
disk[43] <= 32'b001111_11110_01011_0000000000000000; 	// lw
disk[44] <= 32'b000010_01010_11011_0000000000000001; 	// subi
disk[45] <= 32'b010010_11110_11011_1111111111111111; 	// sw
disk[46] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[47] <= 32'b111100_00000000000000000000100100; 	// j
disk[48] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[49] <= 32'b001110_01010_00001_0000000000000000; 	// mov
disk[50] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[51] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[52] <= 32'b010000_00000_10100_0000000000000001; 	// li
disk[53] <= 32'b010010_00101_10100_0000000000000000; 	// sw
disk[54] <= 32'b010000_00000_10101_0000000000000010; 	// li
disk[55] <= 32'b010010_00101_10101_0000000000000001; 	// sw
disk[56] <= 32'b010000_00000_10110_0000000000000011; 	// li
disk[57] <= 32'b010010_00101_10110_0000000000000010; 	// sw
disk[58] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[59] <= 32'b010010_11110_10111_0000000000000000; 	// sw
disk[60] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[61] <= 32'b010000_00000_11001_0000000000001010; 	// li
disk[62] <= 32'b000000_01010_11001_11000_00000_001110; 	// lt
disk[63] <= 32'b010101_11000_00000_0000000001010100; 	// jf
disk[64] <= 32'b010001_00101_01011_0000000000000011; 	// la
disk[65] <= 32'b000000_01011_01010_11010_00000_000000; 	// add
disk[66] <= 32'b010000_00000_11011_0000000000000000; 	// li
disk[67] <= 32'b010010_11010_11011_0000000000000000; 	// sw
disk[68] <= 32'b010001_00101_01100_0000000000001101; 	// la
disk[69] <= 32'b000000_01100_01010_11100_00000_000000; 	// add
disk[70] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[71] <= 32'b010010_11100_11101_0000000000000000; 	// sw
disk[72] <= 32'b010001_00101_01101_0000000000010111; 	// la
disk[73] <= 32'b000000_01101_01010_10100_00000_000000; 	// add
disk[74] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[75] <= 32'b010010_10100_10101_0000000000000000; 	// sw
disk[76] <= 32'b010001_00101_01110_0000000000100001; 	// la
disk[77] <= 32'b000000_01110_01010_10110_00000_000000; 	// add
disk[78] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[79] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[80] <= 32'b000001_01010_11000_0000000000000001; 	// addi
disk[81] <= 32'b010010_11110_11000_0000000000000000; 	// sw
disk[82] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[83] <= 32'b111100_00000000000000000000111100; 	// j
disk[84] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[85] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[86] <= 32'b010000_00000_10100_0000000000100000; 	// li
disk[87] <= 32'b010010_00101_10100_0000000001101100; 	// sw
disk[88] <= 32'b010000_00000_10101_0000000001000000; 	// li
disk[89] <= 32'b010010_00101_10101_0000000001101101; 	// sw
disk[90] <= 32'b010000_00000_10110_0000000001100100; 	// li
disk[91] <= 32'b010010_00101_10110_0000000001101110; 	// sw
disk[92] <= 32'b010000_00000_10111_0000000000001010; 	// li
disk[93] <= 32'b010010_00101_10111_0000000001101111; 	// sw
disk[94] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[95] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[96] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[97] <= 32'b010010_00101_10100_0000000010011101; 	// sw
disk[98] <= 32'b010000_00000_10101_0000000000000001; 	// li
disk[99] <= 32'b010010_00101_10101_0000000010011110; 	// sw
disk[100] <= 32'b010000_00000_10110_0000000000000010; 	// li
disk[101] <= 32'b010010_00101_10110_0000000010011111; 	// sw
disk[102] <= 32'b010000_00000_10111_0000000000000011; 	// li
disk[103] <= 32'b010010_00101_10111_0000000010100000; 	// sw
disk[104] <= 32'b010000_00000_11000_0000000000000100; 	// li
disk[105] <= 32'b010010_00101_11000_0000000010100001; 	// sw
disk[106] <= 32'b010000_00000_11001_0000000000000101; 	// li
disk[107] <= 32'b010010_00101_11001_0000000010100010; 	// sw
disk[108] <= 32'b010000_00000_11010_0000000000001010; 	// li
disk[109] <= 32'b010010_00101_11010_0000000010100011; 	// sw
disk[110] <= 32'b001111_00101_01010_0000000010011101; 	// lw
disk[111] <= 32'b010010_00101_01010_0000000010100100; 	// sw
disk[112] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[113] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[114] <= 32'b010000_00000_10100_0000011111111111; 	// li
disk[115] <= 32'b010010_00101_10100_0000000001110001; 	// sw
disk[116] <= 32'b010000_00000_10101_0000000000011111; 	// li
disk[117] <= 32'b010010_00101_10101_0000000010011010; 	// sw
disk[118] <= 32'b010000_00000_10110_0000000000111101; 	// li
disk[119] <= 32'b010010_00101_10110_0000000010011011; 	// sw
disk[120] <= 32'b010000_00000_10111_0000000000111111; 	// li
disk[121] <= 32'b010010_00101_10111_0000000010011100; 	// sw
disk[122] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[123] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[124] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[125] <= 32'b010010_11110_10100_1111111111111110; 	// sw
disk[126] <= 32'b001111_11110_01010_1111111111111110; 	// lw
disk[127] <= 32'b001111_00101_01011_0000000001101101; 	// lw
disk[128] <= 32'b000000_01010_01011_10101_00000_001110; 	// lt
disk[129] <= 32'b010101_10101_00000_0000000010001010; 	// jf
disk[130] <= 32'b010001_00101_01100_0000000000101100; 	// la
disk[131] <= 32'b000000_01100_01010_10110_00000_000000; 	// add
disk[132] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[133] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[134] <= 32'b000001_01010_11000_0000000000000001; 	// addi
disk[135] <= 32'b010010_11110_11000_1111111111111110; 	// sw
disk[136] <= 32'b001111_11110_01010_1111111111111110; 	// lw
disk[137] <= 32'b111100_00000000000000000001111110; 	// j
disk[138] <= 32'b010010_11110_11111_1111111111111101; 	// sw
disk[139] <= 32'b111110_00000000000000000000000001; 	// jal
disk[140] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[141] <= 32'b001111_11110_11111_1111111111111101; 	// lw
disk[142] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[143] <= 32'b010010_11110_01010_0000000000000000; 	// sw
disk[144] <= 32'b001111_11110_01011_0000000000000000; 	// lw
disk[145] <= 32'b000001_01011_11001_0000000000000001; 	// addi
disk[146] <= 32'b010010_00101_11001_0000000001110000; 	// sw
disk[147] <= 32'b001111_00101_01100_0000000001101100; 	// lw
disk[148] <= 32'b000000_01011_01100_11010_00000_000011; 	// div
disk[149] <= 32'b010010_11110_11010_1111111111111111; 	// sw
disk[150] <= 32'b000000_01011_01100_11011_00000_000100; 	// mod
disk[151] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[152] <= 32'b000000_11011_11101_11100_00000_010000; 	// gt
disk[153] <= 32'b010101_11100_00000_0000000010011110; 	// jf
disk[154] <= 32'b001111_11110_01101_1111111111111111; 	// lw
disk[155] <= 32'b000001_01101_10100_0000000000000001; 	// addi
disk[156] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[157] <= 32'b001111_11110_01101_1111111111111111; 	// lw
disk[158] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[159] <= 32'b010010_11110_10101_1111111111111110; 	// sw
disk[160] <= 32'b001111_11110_01010_1111111111111110; 	// lw
disk[161] <= 32'b001111_11110_01011_1111111111111111; 	// lw
disk[162] <= 32'b000000_01010_01011_10110_00000_001110; 	// lt
disk[163] <= 32'b010101_10110_00000_0000000010101100; 	// jf
disk[164] <= 32'b010001_00101_01100_0000000000101100; 	// la
disk[165] <= 32'b000000_01100_01010_10111_00000_000000; 	// add
disk[166] <= 32'b010000_00000_11000_0000000000000001; 	// li
disk[167] <= 32'b010010_10111_11000_0000000000000000; 	// sw
disk[168] <= 32'b000001_01010_11001_0000000000000001; 	// addi
disk[169] <= 32'b010010_11110_11001_1111111111111110; 	// sw
disk[170] <= 32'b001111_11110_01010_1111111111111110; 	// lw
disk[171] <= 32'b111100_00000000000000000010100000; 	// j
disk[172] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[173] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[174] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[175] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[176] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[177] <= 32'b001111_00101_01011_0000000001101111; 	// lw
disk[178] <= 32'b000000_01010_01011_10101_00000_001110; 	// lt
disk[179] <= 32'b010101_10101_00000_0000000011001000; 	// jf
disk[180] <= 32'b010001_00101_01100_0000000001110010; 	// la
disk[181] <= 32'b000000_01100_01010_10110_00000_000000; 	// add
disk[182] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[183] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[184] <= 32'b010001_00101_01101_0000000001111100; 	// la
disk[185] <= 32'b000000_01101_01010_11000_00000_000000; 	// add
disk[186] <= 32'b010000_00000_11001_0000000000000000; 	// li
disk[187] <= 32'b010010_11000_11001_0000000000000000; 	// sw
disk[188] <= 32'b010001_00101_01110_0000000010000110; 	// la
disk[189] <= 32'b000000_01110_01010_11010_00000_000000; 	// add
disk[190] <= 32'b010000_00000_11011_0000000000000000; 	// li
disk[191] <= 32'b010010_11010_11011_0000000000000000; 	// sw
disk[192] <= 32'b010001_00101_01111_0000000010010000; 	// la
disk[193] <= 32'b000000_01111_01010_11100_00000_000000; 	// add
disk[194] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[195] <= 32'b010010_11100_11101_0000000000000000; 	// sw
disk[196] <= 32'b000001_01010_10100_0000000000000001; 	// addi
disk[197] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[198] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[199] <= 32'b111100_00000000000000000010110000; 	// j
disk[200] <= 32'b001111_00101_01010_0000000001110000; 	// lw
disk[201] <= 32'b010010_11110_01010_1111111111111110; 	// sw
disk[202] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[203] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[204] <= 32'b001111_11110_01010_1111111111111110; 	// lw
disk[205] <= 32'b001111_00101_01011_0000000001110001; 	// lw
disk[206] <= 32'b000000_01010_01011_10110_00000_001110; 	// lt
disk[207] <= 32'b010101_10110_00000_0000000011101000; 	// jf
disk[208] <= 32'b001110_01010_00110_0000000000000000; 	// mov
disk[209] <= 32'b010110_00110_10111_0000000000000000; 	// ldk
disk[210] <= 32'b010010_11110_10111_0000000000000000; 	// sw
disk[211] <= 32'b001111_11110_01100_0000000000000000; 	// lw
disk[212] <= 32'b001101_01100_11000_0000000000011010; 	// srli
disk[213] <= 32'b001111_00101_01101_0000000010011011; 	// lw
disk[214] <= 32'b000000_11000_01101_11001_00000_001100; 	// eq
disk[215] <= 32'b010101_11001_00000_0000000011100011; 	// jf
disk[216] <= 32'b001111_11110_01110_1111111111111111; 	// lw
disk[217] <= 32'b000001_01110_11010_0000000000000001; 	// addi
disk[218] <= 32'b010001_00101_01111_0000000001110010; 	// la
disk[219] <= 32'b000000_01111_01110_11011_00000_000000; 	// add
disk[220] <= 32'b010010_11011_11010_0000000000000000; 	// sw
disk[221] <= 32'b010001_00101_10000_0000000001111100; 	// la
disk[222] <= 32'b000000_10000_01110_11100_00000_000000; 	// add
disk[223] <= 32'b010010_11100_01010_0000000000000000; 	// sw
disk[224] <= 32'b000001_01110_11101_0000000000000001; 	// addi
disk[225] <= 32'b010010_11110_11101_1111111111111111; 	// sw
disk[226] <= 32'b001111_11110_01110_1111111111111111; 	// lw
disk[227] <= 32'b001111_11110_01010_1111111111111110; 	// lw
disk[228] <= 32'b000001_01010_10100_0000000000000001; 	// addi
disk[229] <= 32'b010010_11110_10100_1111111111111110; 	// sw
disk[230] <= 32'b001111_11110_01010_1111111111111110; 	// lw
disk[231] <= 32'b111100_00000000000000000011001100; 	// j
disk[232] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[233] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[234] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[235] <= 32'b111110_00000000000000000000110011; 	// jal
disk[236] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[237] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[238] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[239] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[240] <= 32'b111110_00000000000000000001010101; 	// jal
disk[241] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[242] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[243] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[244] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[245] <= 32'b111110_00000000000000000001011111; 	// jal
disk[246] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[247] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[248] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[249] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[250] <= 32'b111110_00000000000000000001110001; 	// jal
disk[251] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[252] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[253] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[254] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[255] <= 32'b111110_00000000000000000001111011; 	// jal
disk[256] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[257] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[258] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[259] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[260] <= 32'b111110_00000000000000000010101101; 	// jal
disk[261] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[262] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[263] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[264] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[265] <= 32'b000001_11110_11110_0000000000000110; 	// addi
disk[266] <= 32'b010010_11110_00110_1111111111111101; 	// sw
disk[267] <= 32'b001111_11110_01010_1111111111111101; 	// lw
disk[268] <= 32'b001111_00101_01011_0000000001101100; 	// lw
disk[269] <= 32'b000000_01010_01011_10100_00000_000011; 	// div
disk[270] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[271] <= 32'b000000_01010_01011_10101_00000_000100; 	// mod
disk[272] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[273] <= 32'b000000_10101_10111_10110_00000_010000; 	// gt
disk[274] <= 32'b010101_10110_00000_0000000100010111; 	// jf
disk[275] <= 32'b001111_11110_01100_1111111111111111; 	// lw
disk[276] <= 32'b000001_01100_11000_0000000000000001; 	// addi
disk[277] <= 32'b010010_11110_11000_1111111111111111; 	// sw
disk[278] <= 32'b001111_11110_01100_1111111111111111; 	// lw
disk[279] <= 32'b010000_00000_11001_0000000000000000; 	// li
disk[280] <= 32'b010010_11110_11001_1111111111111110; 	// sw
disk[281] <= 32'b001111_11110_01010_1111111111111110; 	// lw
disk[282] <= 32'b001111_00101_01011_0000000001101101; 	// lw
disk[283] <= 32'b000000_01010_01011_11010_00000_001110; 	// lt
disk[284] <= 32'b010101_11010_00000_0000000100111100; 	// jf
disk[285] <= 32'b010001_00101_01100_0000000000101100; 	// la
disk[286] <= 32'b000000_01100_01010_11011_00000_000000; 	// add
disk[287] <= 32'b001111_11011_11011_0000000000000000; 	// lw
disk[288] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[289] <= 32'b000000_11011_11101_11100_00000_001100; 	// eq
disk[290] <= 32'b010101_11100_00000_0000000100110111; 	// jf
disk[291] <= 32'b010010_11110_01010_0000000000000000; 	// sw
disk[292] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[293] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[294] <= 32'b000000_01010_10101_10100_00000_001101; 	// ne
disk[295] <= 32'b010101_10100_00000_0000000100110100; 	// jf
disk[296] <= 32'b010001_00101_01011_0000000000101100; 	// la
disk[297] <= 32'b001111_11110_01100_1111111111111110; 	// lw
disk[298] <= 32'b000000_01011_01100_10110_00000_000000; 	// add
disk[299] <= 32'b010000_00000_10111_0000000000000001; 	// li
disk[300] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[301] <= 32'b000010_01010_11000_0000000000000001; 	// subi
disk[302] <= 32'b010010_11110_11000_1111111111111111; 	// sw
disk[303] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[304] <= 32'b000001_01100_11001_0000000000000001; 	// addi
disk[305] <= 32'b010010_11110_11001_1111111111111110; 	// sw
disk[306] <= 32'b001111_11110_01100_1111111111111110; 	// lw
disk[307] <= 32'b111100_00000000000000000100100100; 	// j
disk[308] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[309] <= 32'b001110_01010_00001_0000000000000000; 	// mov
disk[310] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[311] <= 32'b001111_11110_01010_1111111111111110; 	// lw
disk[312] <= 32'b000001_01010_11010_0000000000000001; 	// addi
disk[313] <= 32'b010010_11110_11010_1111111111111110; 	// sw
disk[314] <= 32'b001111_11110_01010_1111111111111110; 	// lw
disk[315] <= 32'b111100_00000000000000000100011001; 	// j
disk[316] <= 32'b001111_00101_01010_0000000001101110; 	// lw
disk[317] <= 32'b001110_01010_00001_0000000000000000; 	// mov
disk[318] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[319] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[320] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[321] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[322] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[323] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[324] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[325] <= 32'b001111_00101_01011_0000000001101111; 	// lw
disk[326] <= 32'b000000_01010_01011_10110_00000_001110; 	// lt
disk[327] <= 32'b010101_10110_00000_0000000101011101; 	// jf
disk[328] <= 32'b010001_00101_01100_0000000010000110; 	// la
disk[329] <= 32'b000000_01100_01010_10111_00000_000000; 	// add
disk[330] <= 32'b001111_10111_10111_0000000000000000; 	// lw
disk[331] <= 32'b010000_00000_11001_0000000000000000; 	// li
disk[332] <= 32'b000000_10111_11001_11000_00000_001101; 	// ne
disk[333] <= 32'b010101_11000_00000_0000000101011000; 	// jf
disk[334] <= 32'b001110_01010_00110_0000000000000000; 	// mov
disk[335] <= 32'b010010_11110_11111_1111111111111110; 	// sw
disk[336] <= 32'b111110_00000000000000000000011001; 	// jal
disk[337] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[338] <= 32'b001111_11110_11111_1111111111111110; 	// lw
disk[339] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[340] <= 32'b001111_11110_01011_0000000000000000; 	// lw
disk[341] <= 32'b000000_01011_01010_11010_00000_000000; 	// add
disk[342] <= 32'b010010_11110_11010_0000000000000000; 	// sw
disk[343] <= 32'b001111_11110_01011_0000000000000000; 	// lw
disk[344] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[345] <= 32'b000001_01010_11011_0000000000000001; 	// addi
disk[346] <= 32'b010010_11110_11011_1111111111111111; 	// sw
disk[347] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[348] <= 32'b111100_00000000000000000101000100; 	// j
disk[349] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[350] <= 32'b001110_01010_00001_0000000000000000; 	// mov
disk[351] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[352] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[353] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[354] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[355] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[356] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[357] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[358] <= 32'b001111_00101_01011_0000000001101111; 	// lw
disk[359] <= 32'b000000_01010_01011_10110_00000_001110; 	// lt
disk[360] <= 32'b010101_10110_00000_0000000101111110; 	// jf
disk[361] <= 32'b010001_00101_01100_0000000001110010; 	// la
disk[362] <= 32'b000000_01100_01010_10111_00000_000000; 	// add
disk[363] <= 32'b001111_10111_10111_0000000000000000; 	// lw
disk[364] <= 32'b010000_00000_11001_0000000000000000; 	// li
disk[365] <= 32'b000000_10111_11001_11000_00000_001101; 	// ne
disk[366] <= 32'b010101_11000_00000_0000000101111001; 	// jf
disk[367] <= 32'b001110_01010_00110_0000000000000000; 	// mov
disk[368] <= 32'b010010_11110_11111_1111111111111110; 	// sw
disk[369] <= 32'b111110_00000000000000000000011001; 	// jal
disk[370] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[371] <= 32'b001111_11110_11111_1111111111111110; 	// lw
disk[372] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[373] <= 32'b001111_11110_01011_0000000000000000; 	// lw
disk[374] <= 32'b000000_01011_01010_11010_00000_000000; 	// add
disk[375] <= 32'b010010_11110_11010_0000000000000000; 	// sw
disk[376] <= 32'b001111_11110_01011_0000000000000000; 	// lw
disk[377] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[378] <= 32'b000001_01010_11011_0000000000000001; 	// addi
disk[379] <= 32'b010010_11110_11011_1111111111111111; 	// sw
disk[380] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[381] <= 32'b111100_00000000000000000101100101; 	// j
disk[382] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[383] <= 32'b001110_01010_00001_0000000000000000; 	// mov
disk[384] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[385] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[386] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[387] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[388] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[389] <= 32'b001111_00101_01011_0000000001101111; 	// lw
disk[390] <= 32'b000000_01010_01011_10101_00000_001110; 	// lt
disk[391] <= 32'b010101_10101_00000_0000000110010101; 	// jf
disk[392] <= 32'b010001_00101_01100_0000000000000011; 	// la
disk[393] <= 32'b000000_01100_01010_10110_00000_000000; 	// add
disk[394] <= 32'b001111_10110_10110_0000000000000000; 	// lw
disk[395] <= 32'b001111_00101_01101_0000000000000010; 	// lw
disk[396] <= 32'b000000_10110_01101_10111_00000_001100; 	// eq
disk[397] <= 32'b010101_10111_00000_0000000110010000; 	// jf
disk[398] <= 32'b001110_01010_00001_0000000000000000; 	// mov
disk[399] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[400] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[401] <= 32'b000001_01010_11000_0000000000000001; 	// addi
disk[402] <= 32'b010010_11110_11000_0000000000000000; 	// sw
disk[403] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[404] <= 32'b111100_00000000000000000110000100; 	// j
disk[405] <= 32'b001111_00101_01010_0000000001101110; 	// lw
disk[406] <= 32'b001110_01010_00001_0000000000000000; 	// mov
disk[407] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[408] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[409] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[410] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[411] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[412] <= 32'b001111_00101_01011_0000000001101111; 	// lw
disk[413] <= 32'b000000_01010_01011_10101_00000_001110; 	// lt
disk[414] <= 32'b010101_10101_00000_0000000110101100; 	// jf
disk[415] <= 32'b010001_00101_01100_0000000000000011; 	// la
disk[416] <= 32'b000000_01100_01010_10110_00000_000000; 	// add
disk[417] <= 32'b001111_10110_10110_0000000000000000; 	// lw
disk[418] <= 32'b001111_00101_01101_0000000000000001; 	// lw
disk[419] <= 32'b000000_10110_01101_10111_00000_001100; 	// eq
disk[420] <= 32'b010101_10111_00000_0000000110100111; 	// jf
disk[421] <= 32'b001110_01010_00001_0000000000000000; 	// mov
disk[422] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[423] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[424] <= 32'b000001_01010_11000_0000000000000001; 	// addi
disk[425] <= 32'b010010_11110_11000_0000000000000000; 	// sw
disk[426] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[427] <= 32'b111100_00000000000000000110011011; 	// j
disk[428] <= 32'b001111_00101_01010_0000000001101110; 	// lw
disk[429] <= 32'b001110_01010_00001_0000000000000000; 	// mov
disk[430] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[431] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[432] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[433] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[434] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[435] <= 32'b001111_00101_01011_0000000001101111; 	// lw
disk[436] <= 32'b000000_01010_01011_10101_00000_001110; 	// lt
disk[437] <= 32'b010101_10101_00000_0000000111000101; 	// jf
disk[438] <= 32'b010001_00101_01100_0000000010000110; 	// la
disk[439] <= 32'b000000_01100_01010_10110_00000_000000; 	// add
disk[440] <= 32'b001111_10110_10110_0000000000000000; 	// lw
disk[441] <= 32'b010000_00000_11000_0000000000000000; 	// li
disk[442] <= 32'b000000_10110_11000_10111_00000_001101; 	// ne
disk[443] <= 32'b010101_10111_00000_0000000111000000; 	// jf
disk[444] <= 32'b010001_00101_01101_0000000000000011; 	// la
disk[445] <= 32'b000000_01101_01010_11001_00000_000000; 	// add
disk[446] <= 32'b001111_00101_01110_0000000000000001; 	// lw
disk[447] <= 32'b010010_11001_01110_0000000000000000; 	// sw
disk[448] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[449] <= 32'b000001_01010_11010_0000000000000001; 	// addi
disk[450] <= 32'b010010_11110_11010_0000000000000000; 	// sw
disk[451] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[452] <= 32'b111100_00000000000000000110110010; 	// j
disk[453] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[454] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[455] <= 32'b010010_11110_00110_1111111111111110; 	// sw
disk[456] <= 32'b001111_11110_01010_1111111111111110; 	// lw
disk[457] <= 32'b010010_11110_01010_0000000000000000; 	// sw
disk[458] <= 32'b001111_11110_01011_0000000000000000; 	// lw
disk[459] <= 32'b001110_01011_00110_0000000000000000; 	// mov
disk[460] <= 32'b010110_00110_10100_0000000000000000; 	// ldk
disk[461] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[462] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[463] <= 32'b001101_01010_10101_0000000000011010; 	// srli
disk[464] <= 32'b001111_00101_01011_0000000010011010; 	// lw
disk[465] <= 32'b000000_10101_01011_10110_00000_001101; 	// ne
disk[466] <= 32'b010101_10110_00000_0000000111011100; 	// jf
disk[467] <= 32'b001111_11110_01100_0000000000000000; 	// lw
disk[468] <= 32'b000001_01100_10111_0000000000000001; 	// addi
disk[469] <= 32'b010010_11110_10111_0000000000000000; 	// sw
disk[470] <= 32'b001111_11110_01100_0000000000000000; 	// lw
disk[471] <= 32'b001110_01100_00110_0000000000000000; 	// mov
disk[472] <= 32'b010110_00110_11000_0000000000000000; 	// ldk
disk[473] <= 32'b010010_11110_11000_1111111111111111; 	// sw
disk[474] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[475] <= 32'b111100_00000000000000000111001110; 	// j
disk[476] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[477] <= 32'b001111_11110_01011_1111111111111110; 	// lw
disk[478] <= 32'b000000_01010_01011_11001_00000_000001; 	// sub
disk[479] <= 32'b001110_11001_00001_0000000000000000; 	// mov
disk[480] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[481] <= 32'b000001_11110_11110_0000000000001010; 	// addi
disk[482] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[483] <= 32'b001111_11110_01010_1111111111111001; 	// lw
disk[484] <= 32'b000010_01010_10100_0000000000000001; 	// subi
disk[485] <= 32'b010010_11110_10100_1111111111111001; 	// sw
disk[486] <= 32'b001111_11110_01010_1111111111111001; 	// lw
disk[487] <= 32'b010001_00101_01011_0000000001111100; 	// la
disk[488] <= 32'b000000_01011_01010_10101_00000_000000; 	// add
disk[489] <= 32'b001111_10101_10101_0000000000000000; 	// lw
disk[490] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[491] <= 32'b010001_00101_01100_0000000001110010; 	// la
disk[492] <= 32'b000000_01100_01010_10110_00000_000000; 	// add
disk[493] <= 32'b001111_10110_10110_0000000000000000; 	// lw
disk[494] <= 32'b010010_11110_10110_0000000000000000; 	// sw
disk[495] <= 32'b001111_11110_01101_1111111111111111; 	// lw
disk[496] <= 32'b010010_11110_01101_1111111111111010; 	// sw
disk[497] <= 32'b001110_01101_00110_0000000000000000; 	// mov
disk[498] <= 32'b010010_11110_11111_1111111111111000; 	// sw
disk[499] <= 32'b111110_00000000000000000111000110; 	// jal
disk[500] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[501] <= 32'b001111_11110_11111_1111111111111000; 	// lw
disk[502] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[503] <= 32'b010010_11110_01010_1111111111111110; 	// sw
disk[504] <= 32'b001111_11110_01011_1111111111111110; 	// lw
disk[505] <= 32'b001110_01011_00110_0000000000000000; 	// mov
disk[506] <= 32'b010010_11110_11111_1111111111111000; 	// sw
disk[507] <= 32'b111110_00000000000000000100001001; 	// jal
disk[508] <= 32'b000010_11110_11110_0000000000000110; 	// subi
disk[509] <= 32'b001111_11110_11111_1111111111111000; 	// lw
disk[510] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[511] <= 32'b010010_11110_01010_1111111111111101; 	// sw
disk[512] <= 32'b001111_00101_01011_0000000001101100; 	// lw
disk[513] <= 32'b001111_11110_01100_1111111111111101; 	// lw
disk[514] <= 32'b000000_01011_01100_10111_00000_000010; 	// mul
disk[515] <= 32'b010010_11110_10111_1111111111111011; 	// sw
disk[516] <= 32'b001111_11110_01101_1111111111111010; 	// lw
disk[517] <= 32'b001110_01101_00110_0000000000000000; 	// mov
disk[518] <= 32'b010110_00110_11000_0000000000000000; 	// ldk
disk[519] <= 32'b010010_11110_11000_1111111111111100; 	// sw
disk[520] <= 32'b001111_11110_01010_1111111111111100; 	// lw
disk[521] <= 32'b001101_01010_11001_0000000000011010; 	// srli
disk[522] <= 32'b001111_00101_01011_0000000010011010; 	// lw
disk[523] <= 32'b000000_11001_01011_11010_00000_001101; 	// ne
disk[524] <= 32'b010101_11010_00000_0000001000011101; 	// jf
disk[525] <= 32'b001110_01010_00110_0000000000000000; 	// mov
disk[526] <= 32'b001111_11110_01100_1111111111111011; 	// lw
disk[527] <= 32'b001110_01100_00111_0000000000000000; 	// mov
disk[528] <= 32'b011001_00111_00110_0000000000000000; 	// sim
disk[529] <= 32'b001111_11110_01101_1111111111111010; 	// lw
disk[530] <= 32'b000001_01101_11011_0000000000000001; 	// addi
disk[531] <= 32'b010010_11110_11011_1111111111111010; 	// sw
disk[532] <= 32'b001111_11110_01101_1111111111111010; 	// lw
disk[533] <= 32'b001110_01101_00110_0000000000000000; 	// mov
disk[534] <= 32'b010110_00110_11100_0000000000000000; 	// ldk
disk[535] <= 32'b010010_11110_11100_1111111111111100; 	// sw
disk[536] <= 32'b001111_11110_01010_1111111111111100; 	// lw
disk[537] <= 32'b000001_01100_11101_0000000000000001; 	// addi
disk[538] <= 32'b010010_11110_11101_1111111111111011; 	// sw
disk[539] <= 32'b001111_11110_01100_1111111111111011; 	// lw
disk[540] <= 32'b111100_00000000000000001000001000; 	// j
disk[541] <= 32'b001111_11110_01010_1111111111111100; 	// lw
disk[542] <= 32'b001110_01010_00110_0000000000000000; 	// mov
disk[543] <= 32'b001111_11110_01011_1111111111111011; 	// lw
disk[544] <= 32'b001110_01011_00111_0000000000000000; 	// mov
disk[545] <= 32'b011001_00111_00110_0000000000000000; 	// sim
disk[546] <= 32'b001111_11110_01100_0000000000000000; 	// lw
disk[547] <= 32'b001110_01100_00110_0000000000000000; 	// mov
disk[548] <= 32'b011110_00110_00000_0000000000000000; 	// mmuSelect
disk[549] <= 32'b001111_00101_01101_0000000001101100; 	// lw
disk[550] <= 32'b001111_11110_01110_1111111111111101; 	// lw
disk[551] <= 32'b000000_01101_01110_10100_00000_000010; 	// mul
disk[552] <= 32'b001110_10100_00110_0000000000000000; 	// mov
disk[553] <= 32'b011010_00000_00110_0000000000000000; 	// mmuLowerIM
disk[554] <= 32'b010001_00101_01111_0000000010000110; 	// la
disk[555] <= 32'b001111_11110_10000_1111111111111001; 	// lw
disk[556] <= 32'b000000_01111_10000_10101_00000_000000; 	// add
disk[557] <= 32'b010010_10101_01100_0000000000000000; 	// sw
disk[558] <= 32'b010001_00101_10001_0000000010010000; 	// la
disk[559] <= 32'b000000_10001_10000_10110_00000_000000; 	// add
disk[560] <= 32'b001111_11110_10010_1111111111111111; 	// lw
disk[561] <= 32'b010010_10110_10010_0000000000000000; 	// sw
disk[562] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[563] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[564] <= 32'b010010_11110_00110_0000000000000000; 	// sw
disk[565] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[566] <= 32'b001110_01010_00110_0000000000000000; 	// mov
disk[567] <= 32'b100011_00000_00110_0000000000000000; 	// lcdCurr
disk[568] <= 32'b001111_00101_01011_0000000010100011; 	// lw
disk[569] <= 32'b001110_01011_00110_0000000000000000; 	// mov
disk[570] <= 32'b100001_00000_00110_0000000000000000; 	// lcd
disk[571] <= 32'b010001_00101_01100_0000000000000011; 	// la
disk[572] <= 32'b001111_00101_01101_0000000000101011; 	// lw
disk[573] <= 32'b000000_01100_01101_10100_00000_000000; 	// add
disk[574] <= 32'b001111_00101_01110_0000000000000000; 	// lw
disk[575] <= 32'b010010_10100_01110_0000000000000000; 	// sw
disk[576] <= 32'b010001_00101_01111_0000000000001101; 	// la
disk[577] <= 32'b000000_01111_01101_10101_00000_000000; 	// add
disk[578] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[579] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[580] <= 32'b001110_01010_00110_0000000000000000; 	// mov
disk[581] <= 32'b011110_00110_00000_0000000000000000; 	// mmuSelect
disk[582] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[583] <= 32'b100000_00000000000000000000000000; 	// exec
disk[584] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[585] <= 32'b001110_00010_10111_0000000000000000; 	// mov
disk[586] <= 32'b010000_00000_11001_0000000001101111; 	// li
disk[587] <= 32'b000000_10111_11001_11000_00000_001100; 	// eq
disk[588] <= 32'b010101_11000_00000_0000001001010011; 	// jf
disk[589] <= 32'b000000_01100_01101_11010_00000_000000; 	// add
disk[590] <= 32'b001111_00101_10000_0000000000000010; 	// lw
disk[591] <= 32'b010010_11010_10000_0000000000000000; 	// sw
disk[592] <= 32'b001110_00011_11011_0000000000000000; 	// mov
disk[593] <= 32'b000000_01111_01101_11100_00000_000000; 	// add
disk[594] <= 32'b010010_11100_11011_0000000000000000; 	// sw
disk[595] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[596] <= 32'b001110_00000_00101_0000000000000000; 	// mov
disk[597] <= 32'b000001_11110_11110_0000000010100111; 	// addi
disk[598] <= 32'b111110_00000000000000000011101001; 	// jal
disk[599] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[600] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[601] <= 32'b001111_00101_01011_0000000010011101; 	// lw
disk[602] <= 32'b001110_01011_00110_0000000000000000; 	// mov
disk[603] <= 32'b100001_00000_00110_0000000000000000; 	// lcd
disk[604] <= 32'b010000_00000_10100_0000000000000001; 	// li
disk[605] <= 32'b010101_10100_00000_0000001100100110; 	// jf
disk[606] <= 32'b010011_00000_10101_0000000000000000; 	// in
disk[607] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[608] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[609] <= 32'b001110_01010_00110_0000000000000000; 	// mov
disk[610] <= 32'b010000_00000_00111_0000000000000000; 	// li
disk[611] <= 32'b010100_00000_00110_0000000000000000; 	// out
disk[612] <= 32'b001111_00101_01011_0000000010100100; 	// lw
disk[613] <= 32'b001111_00101_01100_0000000010011101; 	// lw
disk[614] <= 32'b000000_01011_01100_10110_00000_001100; 	// eq
disk[615] <= 32'b010101_10110_00000_0000001001110110; 	// jf
disk[616] <= 32'b010000_00000_11000_0000000000000011; 	// li
disk[617] <= 32'b000000_01010_11000_10111_00000_010000; 	// gt
disk[618] <= 32'b010101_10111_00000_0000001001101110; 	// jf
disk[619] <= 32'b010010_11110_01100_0000000000000000; 	// sw
disk[620] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[621] <= 32'b111100_00000000000000001001110101; 	// j
disk[622] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[623] <= 32'b010000_00000_11010_0000000000000001; 	// li
disk[624] <= 32'b000000_01010_11010_11001_00000_001110; 	// lt
disk[625] <= 32'b010101_11001_00000_0000001001110101; 	// jf
disk[626] <= 32'b001111_00101_01011_0000000010011101; 	// lw
disk[627] <= 32'b010010_11110_01011_0000000000000000; 	// sw
disk[628] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[629] <= 32'b111100_00000000000000001100100000; 	// j
disk[630] <= 32'b001111_00101_01010_0000000010100100; 	// lw
disk[631] <= 32'b001111_00101_01011_0000000010011110; 	// lw
disk[632] <= 32'b000000_01010_01011_11011_00000_001100; 	// eq
disk[633] <= 32'b010101_11011_00000_0000001010001010; 	// jf
disk[634] <= 32'b001111_11110_01100_0000000000000000; 	// lw
disk[635] <= 32'b010000_00000_11101_0000000000000011; 	// li
disk[636] <= 32'b000000_01100_11101_11100_00000_010000; 	// gt
disk[637] <= 32'b010101_11100_00000_0000001010000010; 	// jf
disk[638] <= 32'b001111_00101_01101_0000000010011101; 	// lw
disk[639] <= 32'b010010_11110_01101_0000000000000000; 	// sw
disk[640] <= 32'b001111_11110_01100_0000000000000000; 	// lw
disk[641] <= 32'b111100_00000000000000001010001001; 	// j
disk[642] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[643] <= 32'b010000_00000_10101_0000000000000001; 	// li
disk[644] <= 32'b000000_01010_10101_10100_00000_001110; 	// lt
disk[645] <= 32'b010101_10100_00000_0000001010001001; 	// jf
disk[646] <= 32'b001111_00101_01011_0000000010011101; 	// lw
disk[647] <= 32'b010010_11110_01011_0000000000000000; 	// sw
disk[648] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[649] <= 32'b111100_00000000000000001100100000; 	// j
disk[650] <= 32'b001111_00101_01010_0000000010100100; 	// lw
disk[651] <= 32'b001111_00101_01011_0000000010011111; 	// lw
disk[652] <= 32'b000000_01010_01011_10110_00000_001100; 	// eq
disk[653] <= 32'b010101_10110_00000_0000001010101011; 	// jf
disk[654] <= 32'b001111_11110_01100_0000000000000000; 	// lw
disk[655] <= 32'b010000_00000_11000_0000000000000001; 	// li
disk[656] <= 32'b000000_01100_11000_10111_00000_001100; 	// eq
disk[657] <= 32'b010101_10111_00000_0000001010011011; 	// jf
disk[658] <= 32'b001111_00101_01101_0000000010100001; 	// lw
disk[659] <= 32'b010010_11110_01101_0000000000000000; 	// sw
disk[660] <= 32'b001111_11110_01100_0000000000000000; 	// lw
disk[661] <= 32'b111110_00000000000000000101100000; 	// jal
disk[662] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[663] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[664] <= 32'b001110_01010_00110_0000000000000000; 	// mov
disk[665] <= 32'b100010_00000_00110_0000000000000000; 	// lcdPgms
disk[666] <= 32'b111100_00000000000000001010101010; 	// j
disk[667] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[668] <= 32'b010000_00000_11010_0000000000000011; 	// li
disk[669] <= 32'b000000_01010_11010_11001_00000_010000; 	// gt
disk[670] <= 32'b010101_11001_00000_0000001010100011; 	// jf
disk[671] <= 32'b001111_00101_01011_0000000010011101; 	// lw
disk[672] <= 32'b010010_11110_01011_0000000000000000; 	// sw
disk[673] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[674] <= 32'b111100_00000000000000001010101010; 	// j
disk[675] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[676] <= 32'b010000_00000_11100_0000000000000001; 	// li
disk[677] <= 32'b000000_01010_11100_11011_00000_001110; 	// lt
disk[678] <= 32'b010101_11011_00000_0000001010101010; 	// jf
disk[679] <= 32'b001111_00101_01011_0000000010011101; 	// lw
disk[680] <= 32'b010010_11110_01011_0000000000000000; 	// sw
disk[681] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[682] <= 32'b111100_00000000000000001100100000; 	// j
disk[683] <= 32'b001111_00101_01010_0000000010100100; 	// lw
disk[684] <= 32'b001111_00101_01011_0000000010100000; 	// lw
disk[685] <= 32'b000000_01010_01011_11101_00000_001100; 	// eq
disk[686] <= 32'b010101_11101_00000_0000001011111000; 	// jf
disk[687] <= 32'b001111_11110_01100_0000000000000000; 	// lw
disk[688] <= 32'b010000_00000_10101_0000000000000001; 	// li
disk[689] <= 32'b000000_01100_10101_10100_00000_001100; 	// eq
disk[690] <= 32'b010101_10100_00000_0000001011101001; 	// jf
disk[691] <= 32'b111110_00000000000000000110101111; 	// jal
disk[692] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[693] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[694] <= 32'b111110_00000000000000000110011000; 	// jal
disk[695] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[696] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[697] <= 32'b010010_00101_01010_0000000000101011; 	// sw
disk[698] <= 32'b001111_00101_01011_0000000000101011; 	// lw
disk[699] <= 32'b000001_01011_10110_0000000000000001; 	// addi
disk[700] <= 32'b001110_10110_00110_0000000000000000; 	// mov
disk[701] <= 32'b111110_00000000000000001000110011; 	// jal
disk[702] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[703] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[704] <= 32'b111110_00000000000000000110011000; 	// jal
disk[705] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[706] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[707] <= 32'b010010_00101_01010_0000000000101011; 	// sw
disk[708] <= 32'b001111_00101_01011_0000000000101011; 	// lw
disk[709] <= 32'b000001_01011_10111_0000000000000001; 	// addi
disk[710] <= 32'b001110_10111_00110_0000000000000000; 	// mov
disk[711] <= 32'b111110_00000000000000001000110011; 	// jal
disk[712] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[713] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[714] <= 32'b010001_00101_01011_0000000000000011; 	// la
disk[715] <= 32'b001111_00101_01100_0000000000101011; 	// lw
disk[716] <= 32'b000000_01011_01100_11000_00000_000000; 	// add
disk[717] <= 32'b010000_00000_11001_0000000000000000; 	// li
disk[718] <= 32'b010010_11000_11001_0000000000000000; 	// sw
disk[719] <= 32'b111110_00000000000000000110000001; 	// jal
disk[720] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[721] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[722] <= 32'b010010_00101_01010_0000000000101011; 	// sw
disk[723] <= 32'b001111_00101_01011_0000000000101011; 	// lw
disk[724] <= 32'b000001_01011_11010_0000000000000001; 	// addi
disk[725] <= 32'b001110_11010_00110_0000000000000000; 	// mov
disk[726] <= 32'b100011_00000_00110_0000000000000000; 	// lcdCurr
disk[727] <= 32'b001111_00101_01100_0000000010100011; 	// lw
disk[728] <= 32'b001110_01100_00110_0000000000000000; 	// mov
disk[729] <= 32'b100001_00000_00110_0000000000000000; 	// lcd
disk[730] <= 32'b000001_01011_11011_0000000000000001; 	// addi
disk[731] <= 32'b001110_11011_00110_0000000000000000; 	// mov
disk[732] <= 32'b010001_00101_01101_0000000000001101; 	// la
disk[733] <= 32'b000000_01101_01011_11100_00000_000000; 	// add
disk[734] <= 32'b001111_11100_11100_0000000000000000; 	// lw
disk[735] <= 32'b001110_11100_00111_0000000000000000; 	// mov
disk[736] <= 32'b011110_00110_00000_0000000000000000; 	// mmuSelect
disk[737] <= 32'b100101_00111_00000_0000000000000000; 	// execAgain
disk[738] <= 32'b010001_00101_01110_0000000000000011; 	// la
disk[739] <= 32'b000000_01110_01011_11101_00000_000000; 	// add
disk[740] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[741] <= 32'b010010_11101_10100_0000000000000000; 	// sw
disk[742] <= 32'b001111_00101_01111_0000000010011101; 	// lw
disk[743] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[744] <= 32'b111100_00000000000000001011110111; 	// j
disk[745] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[746] <= 32'b010000_00000_10110_0000000000000010; 	// li
disk[747] <= 32'b000000_01010_10110_10101_00000_001100; 	// eq
disk[748] <= 32'b010101_10101_00000_0000001011110101; 	// jf
disk[749] <= 32'b111110_00000000000000000100111111; 	// jal
disk[750] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[751] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[752] <= 32'b001110_01010_00110_0000000000000000; 	// mov
disk[753] <= 32'b100010_00000_00110_0000000000000000; 	// lcdPgms
disk[754] <= 32'b001111_00101_01011_0000000010100010; 	// lw
disk[755] <= 32'b010010_11110_01011_0000000000000000; 	// sw
disk[756] <= 32'b111100_00000000000000001011110111; 	// j
disk[757] <= 32'b001111_00101_01010_0000000010011101; 	// lw
disk[758] <= 32'b010010_11110_01010_0000000000000000; 	// sw
disk[759] <= 32'b111100_00000000000000001100100000; 	// j
disk[760] <= 32'b001111_00101_01010_0000000010100100; 	// lw
disk[761] <= 32'b001111_00101_01011_0000000010100001; 	// lw
disk[762] <= 32'b000000_01010_01011_10111_00000_001100; 	// eq
disk[763] <= 32'b010101_10111_00000_0000001100000111; 	// jf
disk[764] <= 32'b001111_11110_01100_0000000000000000; 	// lw
disk[765] <= 32'b010000_00000_11001_0000000000000000; 	// li
disk[766] <= 32'b000000_01100_11001_11000_00000_010000; 	// gt
disk[767] <= 32'b010101_11000_00000_0000001100000100; 	// jf
disk[768] <= 32'b001110_01100_00110_0000000000000000; 	// mov
disk[769] <= 32'b111110_00000000000000000111100001; 	// jal
disk[770] <= 32'b000010_11110_11110_0000000000001010; 	// subi
disk[771] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[772] <= 32'b001111_00101_01010_0000000010011101; 	// lw
disk[773] <= 32'b010010_11110_01010_0000000000000000; 	// sw
disk[774] <= 32'b111100_00000000000000001100100000; 	// j
disk[775] <= 32'b001111_00101_01010_0000000010100100; 	// lw
disk[776] <= 32'b001111_00101_01011_0000000010100010; 	// lw
disk[777] <= 32'b000000_01010_01011_11010_00000_001100; 	// eq
disk[778] <= 32'b010101_11010_00000_0000001100100000; 	// jf
disk[779] <= 32'b001111_11110_01100_0000000000000000; 	// lw
disk[780] <= 32'b010000_00000_11100_0000000000000000; 	// li
disk[781] <= 32'b000000_01100_11100_11011_00000_010000; 	// gt
disk[782] <= 32'b010101_11011_00000_0000001100011110; 	// jf
disk[783] <= 32'b000010_01100_11101_0000000000000001; 	// subi
disk[784] <= 32'b010010_00101_11101_0000000000101011; 	// sw
disk[785] <= 32'b001110_01100_00110_0000000000000000; 	// mov
disk[786] <= 32'b111110_00000000000000001000110011; 	// jal
disk[787] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[788] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[789] <= 32'b001110_00011_10100_0000000000000000; 	// mov
disk[790] <= 32'b001110_10100_00110_0000000000000000; 	// mov
disk[791] <= 32'b010000_00000_00111_0000000000000010; 	// li
disk[792] <= 32'b010100_00000_00110_0000000000000010; 	// out
disk[793] <= 32'b010001_00101_01011_0000000000000011; 	// la
disk[794] <= 32'b001111_00101_01100_0000000000101011; 	// lw
disk[795] <= 32'b000000_01011_01100_10101_00000_000000; 	// add
disk[796] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[797] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[798] <= 32'b001111_00101_01010_0000000010011101; 	// lw
disk[799] <= 32'b010010_11110_01010_0000000000000000; 	// sw
disk[800] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[801] <= 32'b010010_00101_01010_0000000010100100; 	// sw
disk[802] <= 32'b001111_00101_01011_0000000010100100; 	// lw
disk[803] <= 32'b001110_01011_00110_0000000000000000; 	// mov
disk[804] <= 32'b100001_00000_00110_0000000000000000; 	// lcd
disk[805] <= 32'b111100_00000000000000001001011100; 	// j
disk[806] <= 32'b111111_00000000000000000000000000; 	// halt


		// PROGRAMA 1
		disk[1700] <= 32'b111101_00000000000000000000100011;		// Jump to Main
		disk[1701] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[1702] <= 32'b010010_11110_00110_1111111111111100; 	// sw
		disk[1703] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[1704] <= 32'b010010_11110_10100_1111111111111111; 	// sw
		disk[1705] <= 32'b010000_00000_10101_0000000000000001; 	// li
		disk[1706] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[1707] <= 32'b010000_00000_10110_0000000000000000; 	// li
		disk[1708] <= 32'b010010_11110_10110_1111111111111101; 	// sw
		disk[1709] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[1710] <= 32'b001111_11110_01011_1111111111111100; 	// lw
		disk[1711] <= 32'b000000_01010_01011_10111_00000_001111; 	// let
		disk[1712] <= 32'b010101_10111_00000_0000000000100000; 	// jf
		disk[1713] <= 32'b010000_00000_11001_0000000000000001; 	// li
		disk[1714] <= 32'b000000_01010_11001_11000_00000_001111; 	// let
		disk[1715] <= 32'b010101_11000_00000_0000000000010010; 	// jf
		disk[1716] <= 32'b010010_11110_01010_1111111111111110; 	// sw
		disk[1717] <= 32'b111100_00000000000000000000011011; 	// j
		disk[1718] <= 32'b001111_11110_01010_1111111111111111; 	// lw
		disk[1719] <= 32'b001111_11110_01011_0000000000000000; 	// lw
		disk[1720] <= 32'b000000_01010_01011_11010_00000_000000; 	// add
		disk[1721] <= 32'b010010_11110_11010_1111111111111110; 	// sw
		disk[1722] <= 32'b010010_11110_01011_1111111111111111; 	// sw
		disk[1723] <= 32'b001111_11110_01010_1111111111111111; 	// lw
		disk[1724] <= 32'b001111_11110_01100_1111111111111110; 	// lw
		disk[1725] <= 32'b010010_11110_01100_0000000000000000; 	// sw
		disk[1726] <= 32'b001111_11110_01011_0000000000000000; 	// lw
		disk[1727] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[1728] <= 32'b000001_01010_11011_0000000000000001; 	// addi
		disk[1729] <= 32'b010010_11110_11011_1111111111111101; 	// sw
		disk[1730] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[1731] <= 32'b111100_00000000000000000000001001; 	// j
		disk[1732] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[1733] <= 32'b001110_01010_00001_0000000000000000; 	// mov
		disk[1734] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1735] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[1736] <= 32'b010000_00000_10100_0000000000001011; 	// li
		disk[1737] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[1738] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[1739] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[1740] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1741] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[1742] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[1743] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1744] <= 32'b001110_00001_01010_0000000000000000; 	// mov
		disk[1745] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[1746] <= 32'b010000_00000_00111_0000000000000000; 	// li
		disk[1747] <= 32'b010100_00000_00110_0000000000000000; 	// out
		disk[1748] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[1749] <= 32'b011111_11111_00000_0000000000000000; 	// syscall
		
		// PROGRAMA 2
		disk[1800] <= 32'b111101_00000000000000000000100001;		// Jump to Main
		disk[1801] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[1802] <= 32'b010010_11110_00110_1111111111111100; 	// sw
		disk[1803] <= 32'b010010_11110_00111_1111111111111101; 	// sw
		disk[1804] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[1805] <= 32'b010010_11110_10100_1111111111111110; 	// sw
		disk[1806] <= 32'b010000_00000_10101_0000000000000000; 	// li
		disk[1807] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[1808] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[1809] <= 32'b001111_11110_01011_1111111111111101; 	// lw
		disk[1810] <= 32'b000000_01010_01011_10110_00000_001110; 	// lt
		disk[1811] <= 32'b010101_10110_00000_0000000000011100; 	// jf
		disk[1812] <= 32'b001111_11110_01100_1111111111111100; 	// lw
		disk[1813] <= 32'b000000_01100_01010_10111_00000_000000; 	// add
		disk[1814] <= 32'b001111_10111_10111_0000000000000000; 	// lw
		disk[1815] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[1816] <= 32'b000000_01101_10111_11000_00000_001110; 	// lt
		disk[1817] <= 32'b010101_11000_00000_0000000000010111; 	// jf
		disk[1818] <= 32'b000000_01100_01010_11001_00000_000000; 	// add
		disk[1819] <= 32'b001111_11001_11001_0000000000000000; 	// lw
		disk[1820] <= 32'b010010_11110_11001_0000000000000000; 	// sw
		disk[1821] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[1822] <= 32'b010010_11110_01010_1111111111111111; 	// sw
		disk[1823] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[1824] <= 32'b000001_01010_11010_0000000000000001; 	// addi
		disk[1825] <= 32'b010010_11110_11010_1111111111111110; 	// sw
		disk[1826] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[1827] <= 32'b111100_00000000000000000000001000; 	// j
		disk[1828] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[1829] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[1830] <= 32'b010000_00000_00111_0000000000000001; 	// li
		disk[1831] <= 32'b010100_00000_00110_0000000000000001; 	// out
		disk[1832] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1833] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[1834] <= 32'b010001_11110_01010_1111111111111011; 	// la
		disk[1835] <= 32'b010000_00000_10100_0000000000001100; 	// li
		disk[1836] <= 32'b010010_01010_10100_0000000000000000; 	// sw
		disk[1837] <= 32'b010000_00000_10101_0000000000101001; 	// li
		disk[1838] <= 32'b010010_01010_10101_0000000000000001; 	// sw
		disk[1839] <= 32'b010000_00000_10110_0000000000010111; 	// li
		disk[1840] <= 32'b010010_01010_10110_0000000000000010; 	// sw
		disk[1841] <= 32'b010000_00000_10111_0000000001100010; 	// li
		disk[1842] <= 32'b010010_01010_10111_0000000000000011; 	// sw
		disk[1843] <= 32'b010000_00000_11000_0000000000100001; 	// li
		disk[1844] <= 32'b010010_01010_11000_0000000000000100; 	// sw
		disk[1845] <= 32'b010000_00000_11001_0000000000010101; 	// li
		disk[1846] <= 32'b010010_01010_11001_0000000000000101; 	// sw
		disk[1847] <= 32'b010001_11110_00110_1111111111111011; 	// la
		disk[1848] <= 32'b010000_00000_00111_0000000000000110; 	// li
		disk[1849] <= 32'b010010_11110_11111_1111111111111010; 	// sw
		disk[1850] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[1851] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[1852] <= 32'b001111_11110_11111_1111111111111010; 	// lw
		disk[1853] <= 32'b001110_00001_01010_0000000000000000; 	// mov
		disk[1854] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[1855] <= 32'b011111_11111_00000_0000000000000000; 	// syscall
		
		// PROGRAMA 3
		disk[1900] <= 32'b111101_00000000000000000000010100;		// Jump to Main
		disk[1901] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[1902] <= 32'b010010_11110_00110_1111111111111111; 	// sw
		disk[1903] <= 32'b010000_00000_10100_0000000000000001; 	// li
		disk[1904] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[1905] <= 32'b001111_11110_01010_1111111111111111; 	// lw
		disk[1906] <= 32'b010000_00000_10110_0000000000000000; 	// li
		disk[1907] <= 32'b000000_01010_10110_10101_00000_010000; 	// gt
		disk[1908] <= 32'b010101_10101_00000_0000000000010001; 	// jf
		disk[1909] <= 32'b001111_11110_01011_0000000000000000; 	// lw
		disk[1910] <= 32'b000000_01011_01010_10111_00000_000010; 	// mul
		disk[1911] <= 32'b010010_11110_10111_0000000000000000; 	// sw
		disk[1912] <= 32'b001111_11110_01011_0000000000000000; 	// lw
		disk[1913] <= 32'b000010_01010_11000_0000000000000001; 	// subi
		disk[1914] <= 32'b010010_11110_11000_1111111111111111; 	// sw
		disk[1915] <= 32'b001111_11110_01010_1111111111111111; 	// lw
		disk[1916] <= 32'b111100_00000000000000000000000101; 	// j
		disk[1917] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[1918] <= 32'b001110_01010_00001_0000000000000000; 	// mov
		disk[1919] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1920] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[1921] <= 32'b001110_11110_00100_0000000000000000; 	// mov
		disk[1922] <= 32'b010000_00000_00010_0000000001101111; 	// li
		disk[1923] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[1924] <= 32'b100100_11111_00011_0000000000000000; 	// block
		disk[1925] <= 32'b010011_00000_10100_0000000000000000; 	// in
		disk[1926] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[1927] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[1928] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[1929] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1930] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[1931] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[1932] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1933] <= 32'b001110_00001_01010_0000000000000000; 	// mov
		disk[1934] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[1935] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[1936] <= 32'b010100_00000_00110_0000000000000010; 	// out
		disk[1937] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[1938] <= 32'b011111_11111_00000_0000000000000000; 	// syscall
		
		//prog 1
		disk[1962] <= 32'b111101_00000000000000000000100011;		// Jump to Main
disk[1963] <= 32'b000001_11110_11110_0000000000000111; 	// addi
disk[1964] <= 32'b010010_11110_00110_1111111111111100; 	// sw
disk[1965] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[1966] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[1967] <= 32'b010000_00000_10101_0000000000000001; 	// li
disk[1968] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[1969] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[1970] <= 32'b010010_11110_10110_1111111111111101; 	// sw
disk[1971] <= 32'b001111_11110_01010_1111111111111101; 	// lw
disk[1972] <= 32'b001111_11110_01011_1111111111111100; 	// lw
disk[1973] <= 32'b000000_01010_01011_10111_00000_001111; 	// let
disk[1974] <= 32'b010101_10111_00000_0000000000100000; 	// jf
disk[1975] <= 32'b010000_00000_11001_0000000000000001; 	// li
disk[1976] <= 32'b000000_01010_11001_11000_00000_001111; 	// let
disk[1977] <= 32'b010101_11000_00000_0000000000010010; 	// jf
disk[1978] <= 32'b010010_11110_01010_1111111111111110; 	// sw
disk[1979] <= 32'b111100_00000000000000000000011011; 	// j
disk[1980] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[1981] <= 32'b001111_11110_01011_0000000000000000; 	// lw
disk[1982] <= 32'b000000_01010_01011_11010_00000_000000; 	// add
disk[1983] <= 32'b010010_11110_11010_1111111111111110; 	// sw
disk[1984] <= 32'b010010_11110_01011_1111111111111111; 	// sw
disk[1985] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[1986] <= 32'b001111_11110_01100_1111111111111110; 	// lw
disk[1987] <= 32'b010010_11110_01100_0000000000000000; 	// sw
disk[1988] <= 32'b001111_11110_01011_0000000000000000; 	// lw
disk[1989] <= 32'b001111_11110_01010_1111111111111101; 	// lw
disk[1990] <= 32'b000001_01010_11011_0000000000000001; 	// addi
disk[1991] <= 32'b010010_11110_11011_1111111111111101; 	// sw
disk[1992] <= 32'b001111_11110_01010_1111111111111101; 	// lw
disk[1993] <= 32'b111100_00000000000000000000001001; 	// j
disk[1994] <= 32'b001111_11110_01010_1111111111111110; 	// lw
disk[1995] <= 32'b001110_01010_00001_0000000000000000; 	// mov
disk[1996] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[1997] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[1998] <= 32'b010000_00000_10100_0000000000001011; 	// li
disk[1999] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[2000] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[2001] <= 32'b001110_01010_00110_0000000000000000; 	// mov
disk[2002] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[2003] <= 32'b111110_00000000000000000000000001; 	// jal
disk[2004] <= 32'b000010_11110_11110_0000000000000111; 	// subi
disk[2005] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[2006] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[2007] <= 32'b001110_01010_00110_0000000000000000; 	// mov
disk[2008] <= 32'b010000_00000_00111_0000000000000000; 	// li
disk[2009] <= 32'b010100_00000_00110_0000000000000000; 	// out
disk[2010] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[2011] <= 32'b011111_11111_00000_0000000000000000; 	// syscall


	
		// SORT
		/*disk[1962] <= 32'b111101_00000000000000000000110110;		// Jump to Main
		disk[1963] <= 32'b000001_11110_11110_0000000000001000; 	// addi
		disk[1964] <= 32'b010010_11110_00110_1111111111111011; 	// sw
		disk[1965] <= 32'b010010_11110_00111_1111111111111100; 	// sw
		disk[1966] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[1967] <= 32'b010010_11110_10100_1111111111111101; 	// sw
		disk[1968] <= 32'b001111_11110_01010_1111111111111100; 	// lw
		disk[1969] <= 32'b000010_01010_10101_0000000000000001; 	// subi
		disk[1970] <= 32'b001111_11110_01011_1111111111111101; 	// lw
		disk[1971] <= 32'b000000_01011_10101_10110_00000_001110; 	// lt
		disk[1972] <= 32'b010101_10110_00000_0000000000110101; 	// jf
		disk[1973] <= 32'b010010_11110_01011_1111111111111111; 	// sw
		disk[1974] <= 32'b000001_01011_10111_0000000000000001; 	// addi
		disk[1975] <= 32'b010010_11110_10111_1111111111111110; 	// sw
		disk[1976] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[1977] <= 32'b001111_11110_01011_1111111111111100; 	// lw
		disk[1978] <= 32'b000000_01010_01011_11000_00000_001110; 	// lt
		disk[1979] <= 32'b010101_11000_00000_0000000000100001; 	// jf
		disk[1980] <= 32'b001111_11110_01100_1111111111111011; 	// lw
		disk[1981] <= 32'b000000_01100_01010_11001_00000_000000; 	// add
		disk[1982] <= 32'b001111_11001_11001_0000000000000000; 	// lw
		disk[1983] <= 32'b001111_11110_01101_1111111111111111; 	// lw
		disk[1984] <= 32'b000000_01100_01101_11010_00000_000000; 	// add
		disk[1985] <= 32'b001111_11010_11010_0000000000000000; 	// lw
		disk[1986] <= 32'b000000_11001_11010_11011_00000_001110; 	// lt
		disk[1987] <= 32'b010101_11011_00000_0000000000011100; 	// jf
		disk[1988] <= 32'b010010_11110_01010_1111111111111111; 	// sw
		disk[1989] <= 32'b001111_11110_01101_1111111111111111; 	// lw
		disk[1990] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[1991] <= 32'b000001_01010_11100_0000000000000001; 	// addi
		disk[1992] <= 32'b010010_11110_11100_1111111111111110; 	// sw
		disk[1993] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[1994] <= 32'b111100_00000000000000000000001110; 	// j
		disk[1995] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[1996] <= 32'b001111_11110_01011_1111111111111111; 	// lw
		disk[1997] <= 32'b000000_01010_01011_11101_00000_001101; 	// ne
		disk[1998] <= 32'b010101_11101_00000_0000000000110000; 	// jf
		disk[1999] <= 32'b001111_11110_01100_1111111111111011; 	// lw
		disk[2000] <= 32'b000000_01100_01010_10100_00000_000000; 	// add
		disk[2001] <= 32'b001111_10100_10100_0000000000000000; 	// lw
		disk[2002] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[2003] <= 32'b000000_01100_01011_10101_00000_000000; 	// add
		disk[2004] <= 32'b001111_10101_10101_0000000000000000; 	// lw
		disk[2005] <= 32'b000000_01100_01010_10110_00000_000000; 	// add
		disk[2006] <= 32'b010010_10110_10101_0000000000000000; 	// sw
		disk[2007] <= 32'b000000_01100_01011_10111_00000_000000; 	// add
		disk[2008] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[2009] <= 32'b010010_10111_01101_0000000000000000; 	// sw
		disk[2010] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[2011] <= 32'b000001_01010_11000_0000000000000001; 	// addi
		disk[2012] <= 32'b010010_11110_11000_1111111111111101; 	// sw
		disk[2013] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[2014] <= 32'b111100_00000000000000000000000110; 	// j
		disk[2015] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[2016] <= 32'b000001_11110_11110_0000000000000110; 	// addi
		disk[2017] <= 32'b010001_11110_01010_1111111111111100; 	// la
		disk[2018] <= 32'b010000_00000_10100_0000000000001001; 	// li
		disk[2019] <= 32'b010010_01010_10100_0000000000000000; 	// sw
		disk[2020] <= 32'b010000_00000_10101_0000000000000110; 	// li
		disk[2021] <= 32'b010010_01010_10101_0000000000000001; 	// sw
		disk[2022] <= 32'b010000_00000_10110_0000000000001000; 	// li
		disk[2023] <= 32'b010010_01010_10110_0000000000000010; 	// sw
		disk[2024] <= 32'b010000_00000_10111_0000000000000111; 	// li
		disk[2025] <= 32'b010010_01010_10111_0000000000000011; 	// sw
		disk[2026] <= 32'b010001_11110_00110_1111111111111100; 	// la
		disk[2027] <= 32'b010000_00000_00111_0000000000000100; 	// li
		disk[2028] <= 32'b010010_11110_11111_1111111111111011; 	// sw
		disk[2029] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[2030] <= 32'b000010_11110_11110_0000000000001000; 	// subi
		disk[2031] <= 32'b001111_11110_11111_1111111111111011; 	// lw
		disk[2032] <= 32'b001110_00001_01010_0000000000000000; 	// mov
		disk[2033] <= 32'b001110_11110_00100_0000000000000000; 	// mov
		disk[2034] <= 32'b010000_00000_00010_0000000001101111; 	// li
		disk[2035] <= 32'b000010_11110_11110_0000000000000110; 	// subi
		disk[2036] <= 32'b100100_11111_00000_0000000000000000; 	// block
		disk[2037] <= 32'b010011_00000_10100_0000000000000000; 	// in
		disk[2038] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[2039] <= 32'b010001_11110_01010_1111111111111100; 	// la
		disk[2040] <= 32'b001111_11110_01011_0000000000000000; 	// lw
		disk[2041] <= 32'b000000_01010_01011_10101_00000_000000; 	// add
		disk[2042] <= 32'b001111_10101_10101_0000000000000000; 	// lw
		disk[2043] <= 32'b001110_10101_00110_0000000000000000; 	// mov
		disk[2044] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[2045] <= 32'b010100_00000_00110_0000000000000010; 	// out
		disk[2046] <= 32'b000010_11110_11110_0000000000000110; 	// subi
		disk[2047] <= 32'b011111_11111_00000_0000000000000000; 	// syscall*/

	end
endmodule
