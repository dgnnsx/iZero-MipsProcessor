library verilog;
use verilog.vl_types.all;
entity BCD_dois_digitos_vlg_vec_tst is
end BCD_dois_digitos_vlg_vec_tst;
