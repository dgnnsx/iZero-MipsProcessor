library verilog;
use verilog.vl_types.all;
entity somador_pc_vlg_vec_tst is
end somador_pc_vlg_vec_tst;
