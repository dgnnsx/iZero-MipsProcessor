module disco_rigido (clk, we, addr, datain, dataout);
	input clk;										// clock
	input we;										// write enable
	input [31:0] addr;							// disk address
	input [31:0] datain;							// data in (to disk)
	
	output reg [31:0] dataout;					// data out (from disk)
	
	localparam DISK_SIZE = 500;				// Tamanho do disco
	reg [31:0] disk [DISK_SIZE-1:0];			// disk cells
	
	always @ (posedge clk) begin
		if (we) disk[addr] <= datain;			// write disk
	end
	
	always @ (negedge clk) begin
		dataout <= disk[addr];
	end

	initial begin
		// SISTEMA OPERACIONAL
		disk[0] <= 32'b010110_00000000000000000000101011;		// Jump to Main
disk[1] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[2] <= 32'b010000_00000_00110_0000000000000000; 	// li
disk[3] <= 32'b010000_00000_00111_0000000000000000; 	// li
disk[4] <= 32'b010100_00000_00110_0000000000000000; 	// out
disk[5] <= 32'b010000_00000_00110_0000000000000000; 	// li
disk[6] <= 32'b010000_00000_00111_0000000000000001; 	// li
disk[7] <= 32'b010100_00000_00110_0000000000000001; 	// out
disk[8] <= 32'b010000_00000_00110_0000000000000000; 	// li
disk[9] <= 32'b010000_00000_00111_0000000000000010; 	// li
disk[10] <= 32'b010100_00000_00110_0000000000000010; 	// out
disk[11] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[12] <= 32'b000001_11110_11110_0000000000000110; 	// addi
disk[13] <= 32'b010010_11110_00110_1111111111111101; 	// sw
disk[14] <= 32'b010000_00000_10100_0000000000100010; 	// li
disk[15] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[16] <= 32'b001111_11110_01010_1111111111111101; 	// lw
disk[17] <= 32'b010010_11110_01010_1111111111111111; 	// sw
disk[18] <= 32'b001111_11110_01011_1111111111111111; 	// lw
disk[19] <= 32'b001110_01011_00110_0000000000000000; 	// mov
disk[20] <= 32'b011001_00110_10101_0000000000000000; 	// ldk
disk[21] <= 32'b010010_11110_10101_1111111111111110; 	// sw
disk[22] <= 32'b001111_11110_01100_1111111111111110; 	// lw
disk[23] <= 32'b001101_01100_10110_0000000000011010; 	// srli
disk[24] <= 32'b001111_11110_01101_0000000000000000; 	// lw
disk[25] <= 32'b000000_10110_01101_10111_00000_001101; 	// ne
disk[26] <= 32'b010101_10111_00000_0000000000100110; 	// jf
disk[27] <= 32'b001110_01100_00110_0000000000000000; 	// mov
disk[28] <= 32'b001110_01011_00111_0000000000000000; 	// mov
disk[29] <= 32'b011100_00111_00110_0000000000000000; 	// sim
disk[30] <= 32'b000001_01011_11000_0000000000000001; 	// addi
disk[31] <= 32'b010010_11110_11000_1111111111111111; 	// sw
disk[32] <= 32'b001111_11110_01011_1111111111111111; 	// lw
disk[33] <= 32'b001110_01011_00110_0000000000000000; 	// mov
disk[34] <= 32'b011001_00110_11001_0000000000000000; 	// ldk
disk[35] <= 32'b010010_11110_11001_1111111111111110; 	// sw
disk[36] <= 32'b001111_11110_01100_1111111111111110; 	// lw
disk[37] <= 32'b010110_00000000000000000000010110; 	// j
disk[38] <= 32'b001110_01100_00110_0000000000000000; 	// mov
disk[39] <= 32'b001110_01011_00111_0000000000000000; 	// mov
disk[40] <= 32'b011100_00111_00110_0000000000000000; 	// sim
disk[41] <= 32'b001110_01011_00001_0000000000000000; 	// mov
disk[42] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[43] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[44] <= 32'b010000_00000_10100_0000000001100011; 	// li
disk[45] <= 32'b010010_11110_10100_1111111111111110; 	// sw
disk[46] <= 32'b010000_00000_10101_0000000010111100; 	// li
disk[47] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[48] <= 32'b001111_11110_01010_1111111111111110; 	// lw
disk[49] <= 32'b001110_01010_00110_0000000000000000; 	// mov
disk[50] <= 32'b010010_11110_01010_1111111111111110; 	// sw
disk[51] <= 32'b010111_00000000000000000000001100; 	// jal
disk[52] <= 32'b001110_00001_01011_0000000000000000; 	// mov
disk[53] <= 32'b000010_11110_11110_0000000000000110; 	// subi
disk[54] <= 32'b001111_11110_01010_1111111111111110; 	// lw
disk[55] <= 32'b010010_11110_01011_1111111111111101; 	// sw
disk[56] <= 32'b001111_11110_01100_1111111111111111; 	// lw
disk[57] <= 32'b001110_01100_00110_0000000000000000; 	// mov
disk[58] <= 32'b010010_11110_01010_1111111111111110; 	// sw
disk[59] <= 32'b010010_11110_01011_1111111111111100; 	// sw
disk[60] <= 32'b010010_11110_01100_1111111111111111; 	// sw
disk[61] <= 32'b010111_00000000000000000000001100; 	// jal
disk[62] <= 32'b001110_00001_01101_0000000000000000; 	// mov
disk[63] <= 32'b000010_11110_11110_0000000000000110; 	// subi
disk[64] <= 32'b001111_11110_01010_1111111111111110; 	// lw
disk[65] <= 32'b001111_11110_01011_1111111111111100; 	// lw
disk[66] <= 32'b001111_11110_01100_1111111111111111; 	// lw
disk[67] <= 32'b010010_11110_01101_1111111111111101; 	// sw
disk[68] <= 32'b010011_00000_10110_0000000000000000; 	// in
disk[69] <= 32'b010010_11110_10110_0000000000000000; 	// sw
disk[70] <= 32'b001111_11110_01110_0000000000000000; 	// lw
disk[71] <= 32'b001110_01110_00110_0000000000000000; 	// mov
disk[72] <= 32'b010000_00000_00111_0000000000000001; 	// li
disk[73] <= 32'b100000_00111_00110_0000000000000000; 	// mmuLower
disk[74] <= 32'b001110_01110_00110_0000000000000000; 	// mov
disk[75] <= 32'b010000_00000_00111_0000000000000000; 	// li
disk[76] <= 32'b010100_00000_00110_0000000000000000; 	// out
disk[77] <= 32'b010000_00000_00110_0000000000000000; 	// li
disk[78] <= 32'b000000_00110_00000_00000_00000_010011; 	// exec
disk[79] <= 32'b011000_00000000000000000000000000; 	// halt

		// MAIOR ELEMENTO
		disk[99] <= 32'b010110_00000000000000000000100011;		// Jump to Main
		disk[100] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[101] <= 32'b010010_11110_00110_1111111111111100; 	// sw
		disk[102] <= 32'b010010_11110_00111_1111111111111101; 	// sw
		disk[103] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[104] <= 32'b010010_11110_10100_1111111111111110; 	// sw
		disk[105] <= 32'b010000_00000_10101_0000000000000000; 	// li
		disk[106] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[107] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[108] <= 32'b001111_11110_01011_1111111111111101; 	// lw
		disk[109] <= 32'b000000_01010_01011_10110_00000_001110; 	// lt
		disk[110] <= 32'b010101_10110_00000_0000000000011011; 	// jf
		disk[111] <= 32'b001111_11110_01100_1111111111111100; 	// lw
		disk[112] <= 32'b000000_01100_01010_10111_00000_000000; 	// add
		disk[113] <= 32'b001111_10111_10111_0000000000000000; 	// lw
		disk[114] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[115] <= 32'b000000_01101_10111_11000_00000_001110; 	// lt
		disk[116] <= 32'b010101_11000_00000_0000000000010111; 	// jf
		disk[117] <= 32'b000000_01100_01010_11001_00000_000000; 	// add
		disk[118] <= 32'b001111_11001_11001_0000000000000000; 	// lw
		disk[119] <= 32'b010010_11110_11001_0000000000000000; 	// sw
		disk[120] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[121] <= 32'b010010_11110_01010_1111111111111111; 	// sw
		disk[122] <= 32'b000001_01010_11010_0000000000000001; 	// addi
		disk[123] <= 32'b010010_11110_11010_1111111111111110; 	// sw
		disk[124] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[125] <= 32'b010110_00000000000000000000001000; 	// j
		disk[126] <= 32'b001111_11110_01110_1111111111111111; 	// lw
		disk[127] <= 32'b001110_01110_00110_0000000000000000; 	// mov
		disk[128] <= 32'b010000_00000_00111_0000000000000001; 	// li
		disk[129] <= 32'b010100_00000_00110_0000000000000001; 	// out
		disk[130] <= 32'b001110_01101_00110_0000000000000000; 	// mov
		disk[131] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[132] <= 32'b010100_00000_00110_0000000000000010; 	// out
		disk[133] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[134] <= 32'b000001_11110_11110_0000000000000110; 	// addi
		disk[135] <= 32'b010001_11110_01010_1111111111111011; 	// la
		disk[136] <= 32'b010000_00000_10100_0000000000001100; 	// li
		disk[137] <= 32'b010010_01010_10100_0000000000000000; 	// sw
		disk[138] <= 32'b010000_00000_10101_0000000000101001; 	// li
		disk[139] <= 32'b010010_01010_10101_0000000000000001; 	// sw
		disk[140] <= 32'b010000_00000_10110_0000000000010111; 	// li
		disk[141] <= 32'b010010_01010_10110_0000000000000010; 	// sw
		disk[142] <= 32'b010000_00000_10111_0000000001100010; 	// li
		disk[143] <= 32'b010010_01010_10111_0000000000000011; 	// sw
		disk[144] <= 32'b010000_00000_11000_0000000000100001; 	// li
		disk[145] <= 32'b010010_01010_11000_0000000000000100; 	// sw
		disk[146] <= 32'b010000_00000_11001_0000000000010101; 	// li
		disk[147] <= 32'b010010_01010_11001_0000000000000101; 	// sw
		disk[148] <= 32'b010001_11110_00110_1111111111111011; 	// la
		disk[149] <= 32'b010000_00000_00111_0000000000000110; 	// li
		disk[150] <= 32'b010111_00000000000000000000000001; 	// jal
		disk[151] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[152] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[153] <= 32'b100010_00000000000000000000000000; 	// syscall
		
		// SORT
		disk[188] <= 32'b010110_00000000000000000000110000;		// Jump to Main
		disk[189] <= 32'b000001_11110_11110_0000000000001000; 	// addi
		disk[190] <= 32'b010010_11110_00110_1111111111111011; 	// sw
		disk[191] <= 32'b010010_11110_00111_1111111111111100; 	// sw
		disk[192] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[193] <= 32'b010010_11110_10100_1111111111111101; 	// sw
		disk[194] <= 32'b001111_11110_01010_1111111111111100; 	// lw
		disk[195] <= 32'b000010_01010_10101_0000000000000001; 	// subi
		disk[196] <= 32'b001111_11110_01011_1111111111111101; 	// lw
		disk[197] <= 32'b000000_01011_10101_10110_00000_001110; 	// lt
		disk[198] <= 32'b010101_10110_00000_0000000000101111; 	// jf
		disk[199] <= 32'b010010_11110_01011_1111111111111111; 	// sw
		disk[200] <= 32'b000001_01011_10111_0000000000000001; 	// addi
		disk[201] <= 32'b010010_11110_10111_1111111111111110; 	// sw
		disk[202] <= 32'b001111_11110_01100_1111111111111110; 	// lw
		disk[203] <= 32'b000000_01100_01010_11000_00000_001110; 	// lt
		disk[204] <= 32'b010101_11000_00000_0000000000011111; 	// jf
		disk[205] <= 32'b001111_11110_01101_1111111111111011; 	// lw
		disk[206] <= 32'b000000_01101_01100_11001_00000_000000; 	// add
		disk[207] <= 32'b001111_11001_11001_0000000000000000; 	// lw
		disk[208] <= 32'b001111_11110_01110_1111111111111111; 	// lw
		disk[209] <= 32'b000000_01101_01110_11010_00000_000000; 	// add
		disk[210] <= 32'b001111_11010_11010_0000000000000000; 	// lw
		disk[211] <= 32'b000000_11001_11010_11011_00000_001110; 	// lt
		disk[212] <= 32'b010101_11011_00000_0000000000011011; 	// jf
		disk[213] <= 32'b010010_11110_01100_1111111111111111; 	// sw
		disk[214] <= 32'b001111_11110_01110_1111111111111111; 	// lw
		disk[215] <= 32'b000001_01100_11100_0000000000000001; 	// addi
		disk[216] <= 32'b010010_11110_11100_1111111111111110; 	// sw
		disk[217] <= 32'b001111_11110_01100_1111111111111110; 	// lw
		disk[218] <= 32'b010110_00000000000000000000001110; 	// j
		disk[219] <= 32'b000000_01011_01110_11101_00000_001101; 	// ne
		disk[220] <= 32'b010101_11101_00000_0000000000101011; 	// jf
		disk[221] <= 32'b000000_01101_01011_10100_00000_000000; 	// add
		disk[222] <= 32'b001111_10100_10100_0000000000000000; 	// lw
		disk[223] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[224] <= 32'b000000_01101_01110_10101_00000_000000; 	// add
		disk[225] <= 32'b001111_10101_10101_0000000000000000; 	// lw
		disk[226] <= 32'b000000_01101_01011_10110_00000_000000; 	// add
		disk[227] <= 32'b010010_10110_10101_0000000000000000; 	// sw
		disk[228] <= 32'b000000_01101_01110_10111_00000_000000; 	// add
		disk[229] <= 32'b001111_11110_01111_0000000000000000; 	// lw
		disk[230] <= 32'b010010_10111_01111_0000000000000000; 	// sw
		disk[231] <= 32'b000001_01011_11000_0000000000000001; 	// addi
		disk[232] <= 32'b010010_11110_11000_1111111111111101; 	// sw
		disk[233] <= 32'b001111_11110_01011_1111111111111101; 	// lw
		disk[234] <= 32'b010110_00000000000000000000000110; 	// j
		disk[235] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[236] <= 32'b000001_11110_11110_0000000000000101; 	// addi
		disk[237] <= 32'b010001_11110_01010_1111111111111100; 	// la
		disk[238] <= 32'b010000_00000_10100_0000000000001001; 	// li
		disk[239] <= 32'b010010_01010_10100_0000000000000000; 	// sw
		disk[240] <= 32'b010000_00000_10101_0000000000000110; 	// li
		disk[241] <= 32'b010010_01010_10101_0000000000000001; 	// sw
		disk[242] <= 32'b010000_00000_10110_0000000000001000; 	// li
		disk[243] <= 32'b010010_01010_10110_0000000000000010; 	// sw
		disk[244] <= 32'b010000_00000_10111_0000000000000111; 	// li
		disk[245] <= 32'b010010_01010_10111_0000000000000011; 	// sw
		disk[246] <= 32'b010001_11110_00110_1111111111111100; 	// la
		disk[247] <= 32'b010000_00000_00111_0000000000000100; 	// li
		disk[248] <= 32'b010111_00000000000000000000000001; 	// jal
		disk[249] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[250] <= 32'b000010_11110_11110_0000000000001000; 	// subi
		disk[251] <= 32'b010011_00000_11000_0000000000000000; 	// in
		disk[252] <= 32'b010010_11110_11000_0000000000000000; 	// sw
		disk[253] <= 32'b010001_11110_01100_1111111111111100; 	// la
		disk[254] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[255] <= 32'b000000_01100_01101_11001_00000_000000; 	// add
		disk[256] <= 32'b001111_11001_11001_0000000000000000; 	// lw
		disk[257] <= 32'b001110_11001_00110_0000000000000000; 	// mov
		disk[258] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[259] <= 32'b010100_00000_00110_0000000000000010; 	// out
		disk[260] <= 32'b100010_00000000000000000000000000; 	// syscall
	end
endmodule
