module disco_rigido (clk, we, addr, datain, dataout);
	input clk;										// clock
	input we;										// write enable
	input [31:0] addr;							// disk address
	input [31:0] datain;							// data in (to disk)
	
	output reg [31:0] dataout;					// data out (from disk)
	
	localparam DISK_SIZE = 100;				// Tamanho do disco
	reg [31:0] disk [DISK_SIZE-1:0];			// disk cells
	
	always @ (posedge clk) begin
		if (we) disk[addr] <= datain;			// write disk
	end
	
	always @ (negedge clk) begin
		dataout <= disk[addr];
	end

	initial begin
		disk[0] <= 32'b010110_00000000000000000000100001;		// Jump to Main
		disk[1] <= 32'b000001_11110_11110_0000000000000011; 	// addi
		disk[2] <= 32'b010010_11110_00110_0000000000000000; 	// sw
		disk[3] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[4] <= 32'b010000_00000_10101_0000000000000010; 	// li
		disk[5] <= 32'b000000_01010_10101_10100_00000_001110; 	// lt
		disk[6] <= 32'b010101_10100_00000_0000000000001010; 	// jf
		disk[7] <= 32'b010000_00000_10110_0000000000000001; 	// li
		disk[8] <= 32'b001110_10110_00001_0000000000000000; 	// mov
		disk[9] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[10] <= 32'b000010_01010_10111_0000000000000001; 	// subi
		disk[11] <= 32'b001110_10111_00110_0000000000000000; 	// mov
		disk[12] <= 32'b010010_11110_11111_1111111111111110; 	// sw
		disk[13] <= 32'b010010_11110_01010_0000000000000000; 	// sw
		disk[14] <= 32'b010111_00000000000000000000000001; 	// jal
		disk[15] <= 32'b000010_11110_11110_0000000000000011; 	// subi
		disk[16] <= 32'b001111_11110_11111_1111111111111110; 	// lw
		disk[17] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[18] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[19] <= 32'b000010_01010_11000_0000000000000010; 	// subi
		disk[20] <= 32'b001110_11000_00110_0000000000000000; 	// mov
		disk[21] <= 32'b010010_11110_11111_1111111111111110; 	// sw
		disk[22] <= 32'b010010_11110_01010_0000000000000000; 	// sw
		disk[23] <= 32'b010010_11110_01011_1111111111111111; 	// sw
		disk[24] <= 32'b010111_00000000000000000000000001; 	// jal
		disk[25] <= 32'b000010_11110_11110_0000000000000011; 	// subi
		disk[26] <= 32'b001111_11110_11111_1111111111111110; 	// lw
		disk[27] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[28] <= 32'b001111_11110_01011_1111111111111111; 	// lw
		disk[29] <= 32'b001110_00001_01100_0000000000000000; 	// mov
		disk[30] <= 32'b000000_01011_01100_11001_00000_000000; 	// add
		disk[31] <= 32'b001110_11001_00001_0000000000000000; 	// mov
		disk[32] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[33] <= 32'b000001_11110_11110_0000000000000001; 	// addi
		disk[34] <= 32'b010011_00000_10100_0000000000000000; 	// in
		disk[35] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[36] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[37] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[38] <= 32'b010010_11110_01010_0000000000000000; 	// sw
		disk[39] <= 32'b010111_00000000000000000000000001; 	// jal
		disk[40] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[41] <= 32'b000010_11110_11110_0000000000000011; 	// subi
		disk[42] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[43] <= 32'b001110_01011_00110_0000000000000000; 	// mov
		disk[44] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[45] <= 32'b010100_00000_00110_0000000000000010; 	// out
		disk[46] <= 32'b011000_00000000000000000000000000; 	// halt
	end
endmodule
