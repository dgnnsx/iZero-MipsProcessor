module disco_rigido (clk, we, addr, datain, dataout);
	input clk;										// clock
	input we;										// write enable
	input [31:0] addr;							// disk address
	input [31:0] datain;							// data in (to disk)
	
	output reg [31:0] dataout;					// data out (from disk)
	
	localparam DISK_SIZE = 500;				// Tamanho do disco
	reg [31:0] disk [DISK_SIZE-1:0];			// disk cells
	
	always @ (posedge clk) begin
		if (we) disk[addr] <= datain;			// write disk
	end
	
	always @ (negedge clk) begin
		dataout <= disk[addr];
	end

	initial begin
		// SISTEMA OPERACIONAL
		disk[0] <= 32'b010110_00000000000000000000110100;		// Jump to Main
		disk[1] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[2] <= 32'b010000_00000_00110_0000000000000000; 	// li
		disk[3] <= 32'b010000_00000_00111_0000000000000000; 	// li
		disk[4] <= 32'b010100_00000_00110_0000000000000000; 	// out
		disk[5] <= 32'b010000_00000_00110_0000000000000000; 	// li
		disk[6] <= 32'b010000_00000_00111_0000000000000001; 	// li
		disk[7] <= 32'b010100_00000_00110_0000000000000001; 	// out
		disk[8] <= 32'b010000_00000_00110_0000000000000000; 	// li
		disk[9] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[10] <= 32'b010100_00000_00110_0000000000000010; 	// out
		disk[11] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[12] <= 32'b000001_11110_11110_0000000000001000; 	// addi
		disk[13] <= 32'b010010_11110_00110_1111111111111011; 	// sw
		disk[14] <= 32'b010010_11110_00111_1111111111111100; 	// sw
		disk[15] <= 32'b010000_00000_10100_0000000000100100; 	// li
		disk[16] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[17] <= 32'b001111_11110_01010_1111111111111011; 	// lw
		disk[18] <= 32'b010010_11110_01010_1111111111111110; 	// sw
		disk[19] <= 32'b001111_00101_01011_0000000000000000; 	// lw
		disk[20] <= 32'b001111_11110_01100_1111111111111100; 	// lw
		disk[21] <= 32'b000000_01011_01100_10101_00000_000010; 	// mul
		disk[22] <= 32'b010010_11110_10101_1111111111111111; 	// sw
		disk[23] <= 32'b001111_11110_01101_1111111111111110; 	// lw
		disk[24] <= 32'b001110_01101_00110_0000000000000000; 	// mov
		disk[25] <= 32'b011001_00110_10110_0000000000000000; 	// ldk
		disk[26] <= 32'b010010_11110_10110_1111111111111101; 	// sw
		disk[27] <= 32'b001111_11110_01110_1111111111111101; 	// lw
		disk[28] <= 32'b001101_01110_10111_0000000000011010; 	// srli
		disk[29] <= 32'b001111_11110_01111_0000000000000000; 	// lw
		disk[30] <= 32'b000000_10111_01111_11000_00000_001101; 	// ne
		disk[31] <= 32'b010101_11000_00000_0000000000101111; 	// jf
		disk[32] <= 32'b001110_01110_00110_0000000000000000; 	// mov
		disk[33] <= 32'b001111_11110_10000_1111111111111111; 	// lw
		disk[34] <= 32'b001110_10000_00111_0000000000000000; 	// mov
		disk[35] <= 32'b011100_00111_00110_0000000000000000; 	// sim
		disk[36] <= 32'b000001_01101_11001_0000000000000001; 	// addi
		disk[37] <= 32'b010010_11110_11001_1111111111111110; 	// sw
		disk[38] <= 32'b001111_11110_01101_1111111111111110; 	// lw
		disk[39] <= 32'b001110_01101_00110_0000000000000000; 	// mov
		disk[40] <= 32'b011001_00110_11010_0000000000000000; 	// ldk
		disk[41] <= 32'b010010_11110_11010_1111111111111101; 	// sw
		disk[42] <= 32'b001111_11110_01110_1111111111111101; 	// lw
		disk[43] <= 32'b000001_10000_11011_0000000000000001; 	// addi
		disk[44] <= 32'b010010_11110_11011_1111111111111111; 	// sw
		disk[45] <= 32'b001111_11110_10000_1111111111111111; 	// lw
		disk[46] <= 32'b010110_00000000000000000000011011; 	// j
		disk[47] <= 32'b001110_01110_00110_0000000000000000; 	// mov
		disk[48] <= 32'b001110_10000_00111_0000000000000000; 	// mov
		disk[49] <= 32'b011100_00111_00110_0000000000000000; 	// sim
		disk[50] <= 32'b001110_10000_00001_0000000000000000; 	// mov
		disk[51] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[52] <= 32'b000001_00101_11110_0000000000000001; 	// addi
		disk[53] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[54] <= 32'b010000_00000_10100_0000000000100000; 	// li
		disk[55] <= 32'b010010_00101_10100_0000000000000000; 	// sw
		disk[56] <= 32'b010000_00000_10101_0000000010010110; 	// li
		disk[57] <= 32'b010010_11110_10101_1111111111111101; 	// sw
		disk[58] <= 32'b010000_00000_10110_0000000011001000; 	// li
		disk[59] <= 32'b010010_11110_10110_1111111111111110; 	// sw
		disk[60] <= 32'b010000_00000_10111_0000000011111110; 	// li
		disk[61] <= 32'b010010_11110_10111_1111111111111111; 	// sw
		disk[62] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[63] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[64] <= 32'b010000_00000_00111_0000000000000101; 	// li
		disk[65] <= 32'b010010_11110_11111_1111111111111001; 	// sw
		disk[66] <= 32'b010010_11110_01010_1111111111111101; 	// sw
		disk[67] <= 32'b010111_00000000000000000000001100; 	// jal
		disk[68] <= 32'b000010_11110_11110_0000000000001000; 	// subi
		disk[69] <= 32'b001111_11110_11111_1111111111111001; 	// lw
		disk[70] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[71] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[72] <= 32'b001111_11110_01100_1111111111111110; 	// lw
		disk[73] <= 32'b001110_01100_00110_0000000000000000; 	// mov
		disk[74] <= 32'b010000_00000_00111_0000000000001000; 	// li
		disk[75] <= 32'b010010_11110_11111_1111111111111001; 	// sw
		disk[76] <= 32'b010010_11110_01010_1111111111111101; 	// sw
		disk[77] <= 32'b010010_11110_01011_1111111111111010; 	// sw
		disk[78] <= 32'b010010_11110_01100_1111111111111110; 	// sw
		disk[79] <= 32'b010111_00000000000000000000001100; 	// jal
		disk[80] <= 32'b000010_11110_11110_0000000000001000; 	// subi
		disk[81] <= 32'b001111_11110_11111_1111111111111001; 	// lw
		disk[82] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[83] <= 32'b001111_11110_01011_1111111111111010; 	// lw
		disk[84] <= 32'b001111_11110_01100_1111111111111110; 	// lw
		disk[85] <= 32'b001110_00001_01101_0000000000000000; 	// mov
		disk[86] <= 32'b001111_11110_01110_1111111111111111; 	// lw
		disk[87] <= 32'b001110_01110_00110_0000000000000000; 	// mov
		disk[88] <= 32'b010000_00000_00111_0000000000001011; 	// li
		disk[89] <= 32'b010010_11110_11111_1111111111111001; 	// sw
		disk[90] <= 32'b010010_11110_01010_1111111111111101; 	// sw
		disk[91] <= 32'b010010_11110_01011_1111111111111010; 	// sw
		disk[92] <= 32'b010010_11110_01100_1111111111111110; 	// sw
		disk[93] <= 32'b010010_11110_01101_1111111111111010; 	// sw
		disk[94] <= 32'b010010_11110_01110_1111111111111111; 	// sw
		disk[95] <= 32'b010111_00000000000000000000001100; 	// jal
		disk[96] <= 32'b000010_11110_11110_0000000000001000; 	// subi
		disk[97] <= 32'b001111_11110_11111_1111111111111001; 	// lw
		disk[98] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[99] <= 32'b001111_11110_01011_1111111111111010; 	// lw
		disk[100] <= 32'b001111_11110_01100_1111111111111110; 	// lw
		disk[101] <= 32'b001111_11110_01101_1111111111111010; 	// lw
		disk[102] <= 32'b001111_11110_01110_1111111111111111; 	// lw
		disk[103] <= 32'b001110_00001_01111_0000000000000000; 	// mov
		disk[104] <= 32'b001111_00101_10000_0000000000000000; 	// lw
		disk[105] <= 32'b000011_10000_11000_0000000000000101; 	// muli
		disk[106] <= 32'b001110_11000_00110_0000000000000000; 	// mov
		disk[107] <= 32'b010000_00000_00111_0000000000000001; 	// li
		disk[108] <= 32'b100000_00111_00110_0000000000000000; 	// mmuLowerIM
		disk[109] <= 32'b100101_00000000000000000000000000; 	// exec
		disk[110] <= 32'b000011_10000_11001_0000000000001000; 	// muli
		disk[111] <= 32'b001110_11001_00110_0000000000000000; 	// mov
		disk[112] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[113] <= 32'b100000_00111_00110_0000000000000000; 	// mmuLowerIM
		disk[114] <= 32'b100101_00000000000000000000000000; 	// exec
		disk[115] <= 32'b000011_10000_11010_0000000000001011; 	// muli
		disk[116] <= 32'b001110_11010_00110_0000000000000000; 	// mov
		disk[117] <= 32'b010000_00000_00111_0000000000000011; 	// li
		disk[118] <= 32'b100000_00111_00110_0000000000000000; 	// mmuLowerIM
		disk[119] <= 32'b100101_00000000000000000000000000; 	// exec
		disk[120] <= 32'b011000_00000000000000000000000000; 	// halt

		// PROGRAMA 1
		disk[150] <= 32'b010110_00000000000000000000100001;		// Jump to Main
		disk[151] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[152] <= 32'b010010_11110_00110_1111111111111100; 	// sw
		disk[153] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[154] <= 32'b010010_11110_10100_1111111111111111; 	// sw
		disk[155] <= 32'b010000_00000_10101_0000000000000001; 	// li
		disk[156] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[157] <= 32'b010000_00000_10110_0000000000000000; 	// li
		disk[158] <= 32'b010010_11110_10110_1111111111111101; 	// sw
		disk[159] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[160] <= 32'b001111_11110_01011_1111111111111100; 	// lw
		disk[161] <= 32'b000000_01010_01011_10111_00000_001111; 	// let
		disk[162] <= 32'b010101_10111_00000_0000000000011111; 	// jf
		disk[163] <= 32'b010000_00000_11001_0000000000000001; 	// li
		disk[164] <= 32'b000000_01010_11001_11000_00000_001111; 	// let
		disk[165] <= 32'b010101_11000_00000_0000000000010010; 	// jf
		disk[166] <= 32'b010010_11110_01010_1111111111111110; 	// sw
		disk[167] <= 32'b010110_00000000000000000000011011; 	// j
		disk[168] <= 32'b001111_11110_01100_1111111111111111; 	// lw
		disk[169] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[170] <= 32'b000000_01100_01101_11010_00000_000000; 	// add
		disk[171] <= 32'b010010_11110_11010_1111111111111110; 	// sw
		disk[172] <= 32'b010010_11110_01101_1111111111111111; 	// sw
		disk[173] <= 32'b001111_11110_01100_1111111111111111; 	// lw
		disk[174] <= 32'b001111_11110_01110_1111111111111110; 	// lw
		disk[175] <= 32'b010010_11110_01110_0000000000000000; 	// sw
		disk[176] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[177] <= 32'b000001_01010_11011_0000000000000001; 	// addi
		disk[178] <= 32'b010010_11110_11011_1111111111111101; 	// sw
		disk[179] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[180] <= 32'b010110_00000000000000000000001001; 	// j
		disk[181] <= 32'b001110_01110_00001_0000000000000000; 	// mov
		disk[182] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[183] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[184] <= 32'b010000_00000_10100_0000000000001010; 	// li
		disk[185] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[186] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[187] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[188] <= 32'b010010_11110_11111_1111111111111010; 	// sw
		disk[189] <= 32'b010010_11110_01010_0000000000000000; 	// sw
		disk[190] <= 32'b010111_00000000000000000000000001; 	// jal
		disk[191] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[192] <= 32'b001111_11110_11111_1111111111111010; 	// lw
		disk[193] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[194] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[195] <= 32'b001110_01011_00110_0000000000000000; 	// mov
		disk[196] <= 32'b010000_00000_00111_0000000000000000; 	// li
		disk[197] <= 32'b010100_00000_00110_0000000000000000; 	// out
		disk[198] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[199] <= 32'b100100_11111_00000_0000000000000000; 	// syscall
		
		// PROGRAMA 2
		disk[200] <= 32'b010110_00000000000000000000011111;		// Jump to Main
		disk[201] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[202] <= 32'b010010_11110_00110_1111111111111100; 	// sw
		disk[203] <= 32'b010010_11110_00111_1111111111111101; 	// sw
		disk[204] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[205] <= 32'b010010_11110_10100_1111111111111110; 	// sw
		disk[206] <= 32'b010000_00000_10101_0000000000000000; 	// li
		disk[207] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[208] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[209] <= 32'b001111_11110_01011_1111111111111101; 	// lw
		disk[210] <= 32'b000000_01010_01011_10110_00000_001110; 	// lt
		disk[211] <= 32'b010101_10110_00000_0000000000011011; 	// jf
		disk[212] <= 32'b001111_11110_01100_1111111111111100; 	// lw
		disk[213] <= 32'b000000_01100_01010_10111_00000_000000; 	// add
		disk[214] <= 32'b001111_10111_10111_0000000000000000; 	// lw
		disk[215] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[216] <= 32'b000000_01101_10111_11000_00000_001110; 	// lt
		disk[217] <= 32'b010101_11000_00000_0000000000010111; 	// jf
		disk[218] <= 32'b000000_01100_01010_11001_00000_000000; 	// add
		disk[219] <= 32'b001111_11001_11001_0000000000000000; 	// lw
		disk[220] <= 32'b010010_11110_11001_0000000000000000; 	// sw
		disk[221] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[222] <= 32'b010010_11110_01010_1111111111111111; 	// sw
		disk[223] <= 32'b000001_01010_11010_0000000000000001; 	// addi
		disk[224] <= 32'b010010_11110_11010_1111111111111110; 	// sw
		disk[225] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[226] <= 32'b010110_00000000000000000000001000; 	// j
		disk[227] <= 32'b001110_01101_00110_0000000000000000; 	// mov
		disk[228] <= 32'b010000_00000_00111_0000000000000001; 	// li
		disk[229] <= 32'b010100_00000_00110_0000000000000001; 	// out
		disk[230] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[231] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[232] <= 32'b010001_11110_01010_1111111111111011; 	// la
		disk[233] <= 32'b010000_00000_10100_0000000000001100; 	// li
		disk[234] <= 32'b010010_01010_10100_0000000000000000; 	// sw
		disk[235] <= 32'b010000_00000_10101_0000000000101001; 	// li
		disk[236] <= 32'b010010_01010_10101_0000000000000001; 	// sw
		disk[237] <= 32'b010000_00000_10110_0000000000010111; 	// li
		disk[238] <= 32'b010010_01010_10110_0000000000000010; 	// sw
		disk[239] <= 32'b010000_00000_10111_0000000001100010; 	// li
		disk[240] <= 32'b010010_01010_10111_0000000000000011; 	// sw
		disk[241] <= 32'b010000_00000_11000_0000000000100001; 	// li
		disk[242] <= 32'b010010_01010_11000_0000000000000100; 	// sw
		disk[243] <= 32'b010000_00000_11001_0000000000010101; 	// li
		disk[244] <= 32'b010010_01010_11001_0000000000000101; 	// sw
		disk[245] <= 32'b010001_11110_00110_1111111111111011; 	// la
		disk[246] <= 32'b010000_00000_00111_0000000000000110; 	// li
		disk[247] <= 32'b010010_11110_11111_1111111111111010; 	// sw
		disk[248] <= 32'b010111_00000000000000000000000001; 	// jal
		disk[249] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[250] <= 32'b001111_11110_11111_1111111111111010; 	// lw
		disk[251] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[252] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[253] <= 32'b100100_11111_00000_0000000000000000; 	// syscall
		
		// PROGRAMA 3
		disk[254] <= 32'b010110_00000000000000000000010011;		// Jump to Main
		disk[255] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[256] <= 32'b010010_11110_00110_1111111111111111; 	// sw
		disk[257] <= 32'b010000_00000_10100_0000000000000001; 	// li
		disk[258] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[259] <= 32'b001111_11110_01010_1111111111111111; 	// lw
		disk[260] <= 32'b010000_00000_10110_0000000000000000; 	// li
		disk[261] <= 32'b000000_01010_10110_10101_00000_010000; 	// gt
		disk[262] <= 32'b010101_10101_00000_0000000000010001; 	// jf
		disk[263] <= 32'b001111_11110_01011_0000000000000000; 	// lw
		disk[264] <= 32'b000000_01011_01010_10111_00000_000010; 	// mul
		disk[265] <= 32'b010010_11110_10111_0000000000000000; 	// sw
		disk[266] <= 32'b001111_11110_01011_0000000000000000; 	// lw
		disk[267] <= 32'b000010_01010_11000_0000000000000001; 	// subi
		disk[268] <= 32'b010010_11110_11000_1111111111111111; 	// sw
		disk[269] <= 32'b001111_11110_01010_1111111111111111; 	// lw
		disk[270] <= 32'b010110_00000000000000000000000101; 	// j
		disk[271] <= 32'b001110_01011_00001_0000000000000000; 	// mov
		disk[272] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[273] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[274] <= 32'b010000_00000_10100_0000000000000111; 	// li
		disk[275] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[276] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[277] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[278] <= 32'b010010_11110_11111_1111111111111101; 	// sw
		disk[279] <= 32'b010010_11110_01010_0000000000000000; 	// sw
		disk[280] <= 32'b010111_00000000000000000000000001; 	// jal
		disk[281] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[282] <= 32'b001111_11110_11111_1111111111111101; 	// lw
		disk[283] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[284] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[285] <= 32'b001110_01011_00110_0000000000000000; 	// mov
		disk[286] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[287] <= 32'b010100_00000_00110_0000000000000010; 	// out
		disk[288] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[289] <= 32'b100100_11111_00000_0000000000000000; 	// syscall
		
	end
endmodule
