module disco_rigido (clk, we, addr, datain, dataout);
	input clk;										// clock
	input we;										// write enable
	input [31:0] addr;							// disk address
	input [31:0] datain;							// data in (to disk)
	
	output reg [31:0] dataout;					// data out (from disk)
	
	localparam DISK_SIZE = 2048;				// Tamanho do disco
	reg [31:0] disk [DISK_SIZE-1:0];			// disk cells
	
	always @ (posedge clk) begin
		if (we) disk[addr] <= datain;			// write disk
	end
	
	always @ (negedge clk) begin
		dataout <= disk[addr];
	end

	initial begin
		// SISTEMA OPERACIONAL

disk[0] <= 32'b111100_00000000000000010001011011;		// Jump to Main
disk[1] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[2] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[3] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[4] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[5] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[6] <= 32'b010110_00001_10000_0000000000000000; 	// ldk
disk[7] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[8] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[9] <= 32'b001101_00101_10001_0000000000011010; 	// srli
disk[10] <= 32'b001111_11101_00110_0000000100010111; 	// lw
disk[11] <= 32'b000000_10001_00110_10010_00000_001101; 	// ne
disk[12] <= 32'b010101_10010_00000_0000000000010110; 	// jf
disk[13] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[14] <= 32'b000001_00111_10011_0000000000000001; 	// addi
disk[15] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[16] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[17] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[18] <= 32'b010110_00001_10100_0000000000000000; 	// ldk
disk[19] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[20] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[21] <= 32'b111100_00000000000000000000001000; 	// j
disk[22] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[23] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[24] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[25] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[26] <= 32'b010010_11110_00001_1111111111111111; 	// sw
disk[27] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[28] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[29] <= 32'b000000_00101_10000_01111_00000_001100; 	// eq
disk[30] <= 32'b010101_01111_00000_0000000000100010; 	// jf
disk[31] <= 32'b010000_00000_10001_0000000000000001; 	// li
disk[32] <= 32'b001110_10001_11000_0000000000000000; 	// mov
disk[33] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[34] <= 32'b010000_00000_10010_0000000000000001; 	// li
disk[35] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[36] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[37] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[38] <= 32'b000000_00101_10100_10011_00000_010000; 	// gt
disk[39] <= 32'b010101_10011_00000_0000000000110000; 	// jf
disk[40] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[41] <= 32'b000011_00110_10101_0000000000000010; 	// muli
disk[42] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[43] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[44] <= 32'b000010_00101_10110_0000000000000001; 	// subi
disk[45] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[46] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[47] <= 32'b111100_00000000000000000000100100; 	// j
disk[48] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[49] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[50] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[51] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[52] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[53] <= 32'b010000_00000_00010_0000000000000000; 	// li
disk[54] <= 32'b010100_00000_00001_0000000000000000; 	// out
disk[55] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[56] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[57] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[58] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[59] <= 32'b010000_00000_00010_0000000000000010; 	// li
disk[60] <= 32'b010100_00000_00001_0000000000000010; 	// out
disk[61] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[62] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[63] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[64] <= 32'b010010_11101_01111_0000000011101000; 	// sw
disk[65] <= 32'b010000_00000_10000_0000000000000001; 	// li
disk[66] <= 32'b010010_11101_10000_0000000011101001; 	// sw
disk[67] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[68] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[69] <= 32'b010000_00000_01111_0000000000000001; 	// li
disk[70] <= 32'b010010_11101_01111_0000000000000000; 	// sw
disk[71] <= 32'b010000_00000_10000_0000000000000010; 	// li
disk[72] <= 32'b010010_11101_10000_0000000000000001; 	// sw
disk[73] <= 32'b010000_00000_10001_0000000000000011; 	// li
disk[74] <= 32'b010010_11101_10001_0000000000000010; 	// sw
disk[75] <= 32'b010000_00000_10010_0000000110010100; 	// li
disk[76] <= 32'b010010_11101_10010_0000000000000011; 	// sw
disk[77] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[78] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[79] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[80] <= 32'b010000_00000_10101_0000000000001010; 	// li
disk[81] <= 32'b000000_00101_10101_10100_00000_001110; 	// lt
disk[82] <= 32'b010101_10100_00000_0000000001110111; 	// jf
disk[83] <= 32'b010001_11101_00110_0000000000000100; 	// la
disk[84] <= 32'b000000_00110_00101_10110_00000_000000; 	// add
disk[85] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[86] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[87] <= 32'b010001_11101_00111_0000000000001110; 	// la
disk[88] <= 32'b000000_00111_00101_01111_00000_000000; 	// add
disk[89] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[90] <= 32'b010010_01111_10000_0000000000000000; 	// sw
disk[91] <= 32'b010001_11101_01000_0000000000011000; 	// la
disk[92] <= 32'b000000_01000_00101_10001_00000_000000; 	// add
disk[93] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[94] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[95] <= 32'b010001_11101_01001_0000000000100010; 	// la
disk[96] <= 32'b000000_01001_00101_10011_00000_000000; 	// add
disk[97] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[98] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[99] <= 32'b010001_11101_01010_0000000000101100; 	// la
disk[100] <= 32'b000000_01010_00101_10101_00000_000000; 	// add
disk[101] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[102] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[103] <= 32'b010001_11101_01011_0000000001000000; 	// la
disk[104] <= 32'b000000_01011_00101_10111_00000_000000; 	// add
disk[105] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[106] <= 32'b010010_10111_01111_0000000000000000; 	// sw
disk[107] <= 32'b010001_11101_01100_0000000001001010; 	// la
disk[108] <= 32'b000000_01100_00101_10000_00000_000000; 	// add
disk[109] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[110] <= 32'b010010_10000_10001_0000000000000000; 	// sw
disk[111] <= 32'b010001_11101_01101_0000000001010100; 	// la
disk[112] <= 32'b000000_01101_00101_10010_00000_000000; 	// add
disk[113] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[114] <= 32'b010010_10010_10011_0000000000000000; 	// sw
disk[115] <= 32'b000001_00101_10100_0000000000000001; 	// addi
disk[116] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[117] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[118] <= 32'b111100_00000000000000000001001111; 	// j
disk[119] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[120] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[121] <= 32'b010000_00000_01111_0000000000100000; 	// li
disk[122] <= 32'b010010_11101_01111_0000000010100000; 	// sw
disk[123] <= 32'b010000_00000_10000_0000000001000000; 	// li
disk[124] <= 32'b010010_11101_10000_0000000010100001; 	// sw
disk[125] <= 32'b010000_00000_10001_0000000001100100; 	// li
disk[126] <= 32'b010010_11101_10001_0000000010100010; 	// sw
disk[127] <= 32'b010000_00000_10010_0000000000001010; 	// li
disk[128] <= 32'b010010_11101_10010_0000000010100011; 	// sw
disk[129] <= 32'b010000_00000_10011_0000001111100111; 	// li
disk[130] <= 32'b010010_11101_10011_0000000001011110; 	// sw
disk[131] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[132] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[133] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[134] <= 32'b010010_11101_01111_0000000100011000; 	// sw
disk[135] <= 32'b010000_00000_10000_0000000000000001; 	// li
disk[136] <= 32'b010010_11101_10000_0000000100011001; 	// sw
disk[137] <= 32'b010000_00000_10001_0000000000000010; 	// li
disk[138] <= 32'b010010_11101_10001_0000000100011010; 	// sw
disk[139] <= 32'b010000_00000_10010_0000000000000011; 	// li
disk[140] <= 32'b010010_11101_10010_0000000100011011; 	// sw
disk[141] <= 32'b010000_00000_10011_0000000000000100; 	// li
disk[142] <= 32'b010010_11101_10011_0000000100011100; 	// sw
disk[143] <= 32'b010000_00000_10100_0000000000000101; 	// li
disk[144] <= 32'b010010_11101_10100_0000000100011101; 	// sw
disk[145] <= 32'b010000_00000_10101_0000000000000110; 	// li
disk[146] <= 32'b010010_11101_10101_0000000100011110; 	// sw
disk[147] <= 32'b010000_00000_10110_0000000000000111; 	// li
disk[148] <= 32'b010010_11101_10110_0000000100011111; 	// sw
disk[149] <= 32'b010000_00000_10111_0000000000001000; 	// li
disk[150] <= 32'b010010_11101_10111_0000000100100000; 	// sw
disk[151] <= 32'b010000_00000_01111_0000000000011110; 	// li
disk[152] <= 32'b010010_11101_01111_0000000100100001; 	// sw
disk[153] <= 32'b001111_11101_00101_0000000100011000; 	// lw
disk[154] <= 32'b010010_11101_00101_0000000100100010; 	// sw
disk[155] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[156] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[157] <= 32'b010000_00000_01111_0000011111111111; 	// li
disk[158] <= 32'b010010_11101_01111_0000000010100101; 	// sw
disk[159] <= 32'b010000_00000_10000_0000000000011111; 	// li
disk[160] <= 32'b010010_11101_10000_0000000100010101; 	// sw
disk[161] <= 32'b010000_00000_10001_0000000000111101; 	// li
disk[162] <= 32'b010010_11101_10001_0000000100010110; 	// sw
disk[163] <= 32'b010000_00000_10010_0000000000111111; 	// li
disk[164] <= 32'b010010_11101_10010_0000000100010111; 	// sw
disk[165] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[166] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[167] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[168] <= 32'b010010_11110_01111_1111111111111110; 	// sw
disk[169] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[170] <= 32'b001111_11101_00110_0000000010100001; 	// lw
disk[171] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[172] <= 32'b010101_10000_00000_0000000010111001; 	// jf
disk[173] <= 32'b010001_11101_00111_0000000001100000; 	// la
disk[174] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[175] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[176] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[177] <= 32'b010001_11101_01000_0000000010101000; 	// la
disk[178] <= 32'b000000_01000_00101_10011_00000_000000; 	// add
disk[179] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[180] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[181] <= 32'b000001_00101_10101_0000000000000001; 	// addi
disk[182] <= 32'b010010_11110_10101_1111111111111110; 	// sw
disk[183] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[184] <= 32'b111100_00000000000000000010101001; 	// j
disk[185] <= 32'b010010_11110_11111_1111111111111101; 	// sw
disk[186] <= 32'b111110_00000000000000000000000001; 	// jal
disk[187] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[188] <= 32'b001111_11110_11111_1111111111111101; 	// lw
disk[189] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[190] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[191] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[192] <= 32'b000001_00110_10110_0000000000000001; 	// addi
disk[193] <= 32'b010010_11101_10110_0000000010100100; 	// sw
disk[194] <= 32'b001111_11101_00111_0000000010100000; 	// lw
disk[195] <= 32'b000000_00110_00111_10111_00000_000011; 	// div
disk[196] <= 32'b010010_11110_10111_1111111111111111; 	// sw
disk[197] <= 32'b000000_00110_00111_01111_00000_000100; 	// mod
disk[198] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[199] <= 32'b000000_01111_10001_10000_00000_010000; 	// gt
disk[200] <= 32'b010101_10000_00000_0000000011001101; 	// jf
disk[201] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[202] <= 32'b000001_01000_10010_0000000000000001; 	// addi
disk[203] <= 32'b010010_11110_10010_1111111111111111; 	// sw
disk[204] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[205] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[206] <= 32'b010010_11110_10011_1111111111111110; 	// sw
disk[207] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[208] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[209] <= 32'b000000_00101_00110_10100_00000_001110; 	// lt
disk[210] <= 32'b010101_10100_00000_0000000011011011; 	// jf
disk[211] <= 32'b010001_11101_00111_0000000001100000; 	// la
disk[212] <= 32'b000000_00111_00101_10101_00000_000000; 	// add
disk[213] <= 32'b010000_00000_10110_0000000000000001; 	// li
disk[214] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[215] <= 32'b000001_00101_10111_0000000000000001; 	// addi
disk[216] <= 32'b010010_11110_10111_1111111111111110; 	// sw
disk[217] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[218] <= 32'b111100_00000000000000000011001111; 	// j
disk[219] <= 32'b001110_11110_01111_0000000000000000; 	// mov
disk[220] <= 32'b001111_11101_00101_0000000010100000; 	// lw
disk[221] <= 32'b000000_01111_00101_10000_00000_000011; 	// div
disk[222] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[223] <= 32'b001110_11110_10001_0000000000000000; 	// mov
disk[224] <= 32'b000000_10001_00101_10010_00000_000100; 	// mod
disk[225] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[226] <= 32'b000000_10010_10100_10011_00000_010000; 	// gt
disk[227] <= 32'b010101_10011_00000_0000000011101000; 	// jf
disk[228] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[229] <= 32'b000001_00110_10101_0000000000000001; 	// addi
disk[230] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[231] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[232] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[233] <= 32'b010010_11110_10110_1111111111111110; 	// sw
disk[234] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[235] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[236] <= 32'b000000_00101_00110_10111_00000_001110; 	// lt
disk[237] <= 32'b010101_10111_00000_0000000011110110; 	// jf
disk[238] <= 32'b010001_11101_00111_0000000010101000; 	// la
disk[239] <= 32'b000000_00111_00101_01111_00000_000000; 	// add
disk[240] <= 32'b010000_00000_10000_0000000000000001; 	// li
disk[241] <= 32'b010010_01111_10000_0000000000000000; 	// sw
disk[242] <= 32'b000001_00101_10001_0000000000000001; 	// addi
disk[243] <= 32'b010010_11110_10001_1111111111111110; 	// sw
disk[244] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[245] <= 32'b111100_00000000000000000011101010; 	// j
disk[246] <= 32'b001111_11101_00101_0000000010100001; 	// lw
disk[247] <= 32'b000010_00101_10010_0000000000000001; 	// subi
disk[248] <= 32'b010001_11101_00110_0000000010101000; 	// la
disk[249] <= 32'b000000_00110_10010_10011_00000_000000; 	// add
disk[250] <= 32'b010000_00000_10100_0000000000000001; 	// li
disk[251] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[252] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[253] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[254] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[255] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[256] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[257] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[258] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[259] <= 32'b010101_10000_00000_0000000100011000; 	// jf
disk[260] <= 32'b010001_11101_00111_0000000011101101; 	// la
disk[261] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[262] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[263] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[264] <= 32'b010001_11101_01000_0000000011110111; 	// la
disk[265] <= 32'b000000_01000_00101_10011_00000_000000; 	// add
disk[266] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[267] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[268] <= 32'b010001_11101_01001_0000000100000001; 	// la
disk[269] <= 32'b000000_01001_00101_10101_00000_000000; 	// add
disk[270] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[271] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[272] <= 32'b010001_11101_01010_0000000100001011; 	// la
disk[273] <= 32'b000000_01010_00101_10111_00000_000000; 	// add
disk[274] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[275] <= 32'b010010_10111_01111_0000000000000000; 	// sw
disk[276] <= 32'b000001_00101_10000_0000000000000001; 	// addi
disk[277] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[278] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[279] <= 32'b111100_00000000000000000100000000; 	// j
disk[280] <= 32'b001111_11101_00101_0000000010100100; 	// lw
disk[281] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[282] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[283] <= 32'b010010_11110_10001_1111111111111111; 	// sw
disk[284] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[285] <= 32'b001111_11101_00110_0000000010100101; 	// lw
disk[286] <= 32'b000000_00101_00110_10010_00000_001110; 	// lt
disk[287] <= 32'b010101_10010_00000_0000000100111000; 	// jf
disk[288] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[289] <= 32'b010110_00001_10011_0000000000000000; 	// ldk
disk[290] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[291] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[292] <= 32'b001101_00111_10100_0000000000011010; 	// srli
disk[293] <= 32'b001111_11101_01000_0000000100010110; 	// lw
disk[294] <= 32'b000000_10100_01000_10101_00000_001100; 	// eq
disk[295] <= 32'b010101_10101_00000_0000000100110011; 	// jf
disk[296] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[297] <= 32'b000001_01001_10110_0000000000000001; 	// addi
disk[298] <= 32'b010001_11101_01010_0000000011101101; 	// la
disk[299] <= 32'b000000_01010_01001_10111_00000_000000; 	// add
disk[300] <= 32'b010010_10111_10110_0000000000000000; 	// sw
disk[301] <= 32'b010001_11101_01011_0000000011110111; 	// la
disk[302] <= 32'b000000_01011_01001_01111_00000_000000; 	// add
disk[303] <= 32'b010010_01111_00101_0000000000000000; 	// sw
disk[304] <= 32'b000001_01001_10000_0000000000000001; 	// addi
disk[305] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[306] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[307] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[308] <= 32'b000001_00101_10001_0000000000000001; 	// addi
disk[309] <= 32'b010010_11110_10001_1111111111111110; 	// sw
disk[310] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[311] <= 32'b111100_00000000000000000100011100; 	// j
disk[312] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[313] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[314] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[315] <= 32'b111110_00000000000000000001000100; 	// jal
disk[316] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[317] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[318] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[319] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[320] <= 32'b111110_00000000000000000001111000; 	// jal
disk[321] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[322] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[323] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[324] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[325] <= 32'b111110_00000000000000000010000100; 	// jal
disk[326] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[327] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[328] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[329] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[330] <= 32'b111110_00000000000000000010011100; 	// jal
disk[331] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[332] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[333] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[334] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[335] <= 32'b111110_00000000000000000010100110; 	// jal
disk[336] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[337] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[338] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[339] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[340] <= 32'b111110_00000000000000000011111101; 	// jal
disk[341] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[342] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[343] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[344] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[345] <= 32'b000001_11110_11110_0000000000000110; 	// addi
disk[346] <= 32'b010010_11110_00001_1111111111111101; 	// sw
disk[347] <= 32'b001111_11110_00101_1111111111111101; 	// lw
disk[348] <= 32'b001111_11101_00110_0000000010100000; 	// lw
disk[349] <= 32'b000000_00101_00110_01111_00000_000011; 	// div
disk[350] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[351] <= 32'b000000_00101_00110_10000_00000_000100; 	// mod
disk[352] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[353] <= 32'b000000_10000_10010_10001_00000_010000; 	// gt
disk[354] <= 32'b010101_10001_00000_0000000101100111; 	// jf
disk[355] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[356] <= 32'b000001_00111_10011_0000000000000001; 	// addi
disk[357] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[358] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[359] <= 32'b010001_11101_00101_0000000001001010; 	// la
disk[360] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[361] <= 32'b000000_00101_00110_10100_00000_000000; 	// add
disk[362] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[363] <= 32'b010010_10100_00111_0000000000000000; 	// sw
disk[364] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[365] <= 32'b010010_11110_10101_1111111111111110; 	// sw
disk[366] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[367] <= 32'b001111_11101_00110_0000000010100001; 	// lw
disk[368] <= 32'b000000_00101_00110_10110_00000_001110; 	// lt
disk[369] <= 32'b010101_10110_00000_0000000110010001; 	// jf
disk[370] <= 32'b010001_11101_00111_0000000001100000; 	// la
disk[371] <= 32'b000000_00111_00101_10111_00000_000000; 	// add
disk[372] <= 32'b001111_10111_10111_0000000000000000; 	// lw
disk[373] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[374] <= 32'b000000_10111_10000_01111_00000_001100; 	// eq
disk[375] <= 32'b010101_01111_00000_0000000110001100; 	// jf
disk[376] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[377] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[378] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[379] <= 32'b000000_00101_10010_10001_00000_010000; 	// gt
disk[380] <= 32'b010101_10001_00000_0000000110001001; 	// jf
disk[381] <= 32'b010001_11101_00110_0000000001100000; 	// la
disk[382] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[383] <= 32'b000000_00110_00111_10011_00000_000000; 	// add
disk[384] <= 32'b010000_00000_10100_0000000000000001; 	// li
disk[385] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[386] <= 32'b000010_00101_10101_0000000000000001; 	// subi
disk[387] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[388] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[389] <= 32'b000001_00111_10110_0000000000000001; 	// addi
disk[390] <= 32'b010010_11110_10110_1111111111111110; 	// sw
disk[391] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[392] <= 32'b111100_00000000000000000101111001; 	// j
disk[393] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[394] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[395] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[396] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[397] <= 32'b000001_00101_10111_0000000000000001; 	// addi
disk[398] <= 32'b010010_11110_10111_1111111111111110; 	// sw
disk[399] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[400] <= 32'b111100_00000000000000000101101110; 	// j
disk[401] <= 32'b001111_11101_00101_0000000010100010; 	// lw
disk[402] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[403] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[404] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[405] <= 32'b010001_11101_00101_0000000000011000; 	// la
disk[406] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[407] <= 32'b000000_00101_00110_01111_00000_000000; 	// add
disk[408] <= 32'b001111_01111_01111_0000000000000000; 	// lw
disk[409] <= 32'b001111_11101_00111_0000000010100000; 	// lw
disk[410] <= 32'b000000_01111_00111_10000_00000_000011; 	// div
disk[411] <= 32'b000001_10000_10001_0000000000000001; 	// addi
disk[412] <= 32'b010010_11110_10001_1111111111111111; 	// sw
disk[413] <= 32'b000000_00101_00110_10010_00000_000000; 	// add
disk[414] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[415] <= 32'b000000_10010_00111_10011_00000_000100; 	// mod
disk[416] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[417] <= 32'b000000_10011_10101_10100_00000_010000; 	// gt
disk[418] <= 32'b010101_10100_00000_0000000110100111; 	// jf
disk[419] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[420] <= 32'b000001_01000_10110_0000000000000001; 	// addi
disk[421] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[422] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[423] <= 32'b001111_11101_00101_0000000010100001; 	// lw
disk[424] <= 32'b000010_00101_10111_0000000000000001; 	// subi
disk[425] <= 32'b010010_11110_10111_1111111111111110; 	// sw
disk[426] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[427] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[428] <= 32'b000000_00101_10000_01111_00000_010000; 	// gt
disk[429] <= 32'b010101_01111_00000_0000000111001101; 	// jf
disk[430] <= 32'b010001_11101_00110_0000000010101000; 	// la
disk[431] <= 32'b000000_00110_00101_10001_00000_000000; 	// add
disk[432] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[433] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[434] <= 32'b000000_10001_10011_10010_00000_001100; 	// eq
disk[435] <= 32'b010101_10010_00000_0000000111001000; 	// jf
disk[436] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[437] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[438] <= 32'b000000_00101_10101_10100_00000_010000; 	// gt
disk[439] <= 32'b010101_10100_00000_0000000111000101; 	// jf
disk[440] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[441] <= 32'b010010_11110_00110_0000000000000000; 	// sw
disk[442] <= 32'b010001_11101_00111_0000000010101000; 	// la
disk[443] <= 32'b000000_00111_00110_10110_00000_000000; 	// add
disk[444] <= 32'b010000_00000_10111_0000000000000001; 	// li
disk[445] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[446] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[447] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[448] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[449] <= 32'b000010_00110_10000_0000000000000001; 	// subi
disk[450] <= 32'b010010_11110_10000_1111111111111110; 	// sw
disk[451] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[452] <= 32'b111100_00000000000000000110110100; 	// j
disk[453] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[454] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[455] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[456] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[457] <= 32'b000010_00101_10001_0000000000000001; 	// subi
disk[458] <= 32'b010010_11110_10001_1111111111111110; 	// sw
disk[459] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[460] <= 32'b111100_00000000000000000110101010; 	// j
disk[461] <= 32'b001111_11101_00101_0000000010100010; 	// lw
disk[462] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[463] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[464] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[465] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[466] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[467] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[468] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[469] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[470] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[471] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[472] <= 32'b010101_10001_00000_0000000111101110; 	// jf
disk[473] <= 32'b010001_11101_00111_0000000100000001; 	// la
disk[474] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
disk[475] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[476] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[477] <= 32'b000000_10010_10100_10011_00000_001101; 	// ne
disk[478] <= 32'b010101_10011_00000_0000000111101001; 	// jf
disk[479] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[480] <= 32'b010010_11110_11111_1111111111111110; 	// sw
disk[481] <= 32'b111110_00000000000000000000011001; 	// jal
disk[482] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[483] <= 32'b001111_11110_11111_1111111111111110; 	// lw
disk[484] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[485] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[486] <= 32'b000000_00110_00101_10101_00000_000000; 	// add
disk[487] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[488] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[489] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[490] <= 32'b000001_00101_10110_0000000000000001; 	// addi
disk[491] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[492] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[493] <= 32'b111100_00000000000000000111010101; 	// j
disk[494] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[495] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[496] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[497] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[498] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[499] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[500] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[501] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[502] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[503] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[504] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[505] <= 32'b010101_10001_00000_0000001000001111; 	// jf
disk[506] <= 32'b010001_11101_00111_0000000011101101; 	// la
disk[507] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
disk[508] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[509] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[510] <= 32'b000000_10010_10100_10011_00000_001101; 	// ne
disk[511] <= 32'b010101_10011_00000_0000001000001010; 	// jf
disk[512] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[513] <= 32'b010010_11110_11111_1111111111111110; 	// sw
disk[514] <= 32'b111110_00000000000000000000011001; 	// jal
disk[515] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[516] <= 32'b001111_11110_11111_1111111111111110; 	// lw
disk[517] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[518] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[519] <= 32'b000000_00110_00101_10101_00000_000000; 	// add
disk[520] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[521] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[522] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[523] <= 32'b000001_00101_10110_0000000000000001; 	// addi
disk[524] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[525] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[526] <= 32'b111100_00000000000000000111110110; 	// j
disk[527] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[528] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[529] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[530] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[531] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[532] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[533] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[534] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[535] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[536] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[537] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[538] <= 32'b010101_10001_00000_0000001000110000; 	// jf
disk[539] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[540] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
disk[541] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[542] <= 32'b001111_11101_01000_0000000000000010; 	// lw
disk[543] <= 32'b000000_10010_01000_10011_00000_001100; 	// eq
disk[544] <= 32'b010101_10011_00000_0000001000101011; 	// jf
disk[545] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[546] <= 32'b010010_11110_11111_1111111111111110; 	// sw
disk[547] <= 32'b111110_00000000000000000000011001; 	// jal
disk[548] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[549] <= 32'b001111_11110_11111_1111111111111110; 	// lw
disk[550] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[551] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[552] <= 32'b000000_00110_00101_10100_00000_000000; 	// add
disk[553] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[554] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[555] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[556] <= 32'b000001_00101_10101_0000000000000001; 	// addi
disk[557] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[558] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[559] <= 32'b111100_00000000000000001000010111; 	// j
disk[560] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[561] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[562] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[563] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[564] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[565] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[566] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[567] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[568] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[569] <= 32'b010101_10000_00000_0000001001000111; 	// jf
disk[570] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[571] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[572] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[573] <= 32'b001111_11101_01000_0000000000000010; 	// lw
disk[574] <= 32'b000000_10001_01000_10010_00000_001100; 	// eq
disk[575] <= 32'b010101_10010_00000_0000001001000010; 	// jf
disk[576] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[577] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[578] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[579] <= 32'b000001_00101_10011_0000000000000001; 	// addi
disk[580] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[581] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[582] <= 32'b111100_00000000000000001000110110; 	// j
disk[583] <= 32'b001111_11101_00101_0000000000000011; 	// lw
disk[584] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[585] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[586] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[587] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[588] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[589] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[590] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[591] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[592] <= 32'b010101_10000_00000_0000001001011110; 	// jf
disk[593] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[594] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[595] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[596] <= 32'b001111_11101_01000_0000000000000001; 	// lw
disk[597] <= 32'b000000_10001_01000_10010_00000_001100; 	// eq
disk[598] <= 32'b010101_10010_00000_0000001001011001; 	// jf
disk[599] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[600] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[601] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[602] <= 32'b000001_00101_10011_0000000000000001; 	// addi
disk[603] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[604] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[605] <= 32'b111100_00000000000000001001001101; 	// j
disk[606] <= 32'b001111_11101_00101_0000000000000011; 	// lw
disk[607] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[608] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[609] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[610] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[611] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[612] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[613] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[614] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[615] <= 32'b010101_10000_00000_0000001001110111; 	// jf
disk[616] <= 32'b010001_11101_00111_0000000100000001; 	// la
disk[617] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[618] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[619] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[620] <= 32'b000000_10001_10011_10010_00000_001101; 	// ne
disk[621] <= 32'b010101_10010_00000_0000001001110010; 	// jf
disk[622] <= 32'b010001_11101_01000_0000000000000100; 	// la
disk[623] <= 32'b000000_01000_00101_10100_00000_000000; 	// add
disk[624] <= 32'b001111_11101_01001_0000000000000001; 	// lw
disk[625] <= 32'b010010_10100_01001_0000000000000000; 	// sw
disk[626] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[627] <= 32'b000001_00101_10101_0000000000000001; 	// addi
disk[628] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[629] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[630] <= 32'b111100_00000000000000001001100100; 	// j
disk[631] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[632] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[633] <= 32'b010010_11110_00001_1111111111111110; 	// sw
disk[634] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[635] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[636] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[637] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[638] <= 32'b010110_00001_01111_0000000000000000; 	// ldk
disk[639] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[640] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[641] <= 32'b001101_00101_10000_0000000000011010; 	// srli
disk[642] <= 32'b001111_11101_00110_0000000100010101; 	// lw
disk[643] <= 32'b000000_10000_00110_10001_00000_001101; 	// ne
disk[644] <= 32'b010101_10001_00000_0000001010001110; 	// jf
disk[645] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[646] <= 32'b000001_00111_10010_0000000000000001; 	// addi
disk[647] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[648] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[649] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[650] <= 32'b010110_00001_10011_0000000000000000; 	// ldk
disk[651] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[652] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[653] <= 32'b111100_00000000000000001010000000; 	// j
disk[654] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[655] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[656] <= 32'b000000_00101_00110_10100_00000_000001; 	// sub
disk[657] <= 32'b001110_10100_11000_0000000000000000; 	// mov
disk[658] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[659] <= 32'b000001_11110_11110_0000000000001010; 	// addi
disk[660] <= 32'b010010_11110_00001_1111111111111001; 	// sw
disk[661] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[662] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[663] <= 32'b010010_11110_01111_1111111111111001; 	// sw
disk[664] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[665] <= 32'b010010_11101_00101_0000000001011111; 	// sw
disk[666] <= 32'b010001_11101_00110_0000000011110111; 	// la
disk[667] <= 32'b000000_00110_00101_10000_00000_000000; 	// add
disk[668] <= 32'b001111_10000_10000_0000000000000000; 	// lw
disk[669] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[670] <= 32'b010001_11101_00111_0000000011101101; 	// la
disk[671] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[672] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[673] <= 32'b010010_11110_10001_0000000000000000; 	// sw
disk[674] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[675] <= 32'b010010_11110_01000_1111111111111010; 	// sw
disk[676] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[677] <= 32'b010010_11110_11111_1111111111111000; 	// sw
disk[678] <= 32'b111110_00000000000000001001111000; 	// jal
disk[679] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[680] <= 32'b001111_11110_11111_1111111111111000; 	// lw
disk[681] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[682] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[683] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[684] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[685] <= 32'b010010_11110_11111_1111111111111000; 	// sw
disk[686] <= 32'b111110_00000000000000000101011001; 	// jal
disk[687] <= 32'b000010_11110_11110_0000000000000110; 	// subi
disk[688] <= 32'b001111_11110_11111_1111111111111000; 	// lw
disk[689] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[690] <= 32'b010010_11110_00101_1111111111111101; 	// sw
disk[691] <= 32'b010001_11101_00110_0000000000110110; 	// la
disk[692] <= 32'b001111_11101_00111_0000000001011111; 	// lw
disk[693] <= 32'b000000_00110_00111_10010_00000_000000; 	// add
disk[694] <= 32'b001111_11110_01000_1111111111111101; 	// lw
disk[695] <= 32'b010010_10010_01000_0000000000000000; 	// sw
disk[696] <= 32'b001111_11101_01001_0000000010100000; 	// lw
disk[697] <= 32'b000000_01001_01000_10011_00000_000010; 	// mul
disk[698] <= 32'b010010_11110_10011_1111111111111011; 	// sw
disk[699] <= 32'b001111_11110_01010_1111111111111010; 	// lw
disk[700] <= 32'b001110_01010_00001_0000000000000000; 	// mov
disk[701] <= 32'b010110_00001_10100_0000000000000000; 	// ldk
disk[702] <= 32'b010010_11110_10100_1111111111111100; 	// sw
disk[703] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[704] <= 32'b001101_00101_10101_0000000000011010; 	// srli
disk[705] <= 32'b001111_11101_00110_0000000100010101; 	// lw
disk[706] <= 32'b000000_10101_00110_10110_00000_001101; 	// ne
disk[707] <= 32'b010101_10110_00000_0000001011010100; 	// jf
disk[708] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[709] <= 32'b001111_11110_00111_1111111111111011; 	// lw
disk[710] <= 32'b001110_00111_00010_0000000000000000; 	// mov
disk[711] <= 32'b011001_00010_00001_0000000000000000; 	// sim
disk[712] <= 32'b001111_11110_01000_1111111111111010; 	// lw
disk[713] <= 32'b000001_01000_10111_0000000000000001; 	// addi
disk[714] <= 32'b010010_11110_10111_1111111111111010; 	// sw
disk[715] <= 32'b001111_11110_01000_1111111111111010; 	// lw
disk[716] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[717] <= 32'b010110_00001_01111_0000000000000000; 	// ldk
disk[718] <= 32'b010010_11110_01111_1111111111111100; 	// sw
disk[719] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[720] <= 32'b000001_00111_10000_0000000000000001; 	// addi
disk[721] <= 32'b010010_11110_10000_1111111111111011; 	// sw
disk[722] <= 32'b001111_11110_00111_1111111111111011; 	// lw
disk[723] <= 32'b111100_00000000000000001010111111; 	// j
disk[724] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[725] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[726] <= 32'b001111_11110_00110_1111111111111011; 	// lw
disk[727] <= 32'b001110_00110_00010_0000000000000000; 	// mov
disk[728] <= 32'b011001_00010_00001_0000000000000000; 	// sim
disk[729] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[730] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[731] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
disk[732] <= 32'b001111_11101_01000_0000000010100000; 	// lw
disk[733] <= 32'b001111_11110_01001_1111111111111101; 	// lw
disk[734] <= 32'b000000_01000_01001_10001_00000_000010; 	// mul
disk[735] <= 32'b001110_10001_00001_0000000000000000; 	// mov
disk[736] <= 32'b011010_00000_00001_0000000000000000; 	// mmuLowerIM
disk[737] <= 32'b010001_11101_01010_0000000100000001; 	// la
disk[738] <= 32'b001111_11110_01011_1111111111111001; 	// lw
disk[739] <= 32'b000000_01010_01011_10010_00000_000000; 	// add
disk[740] <= 32'b010010_10010_00111_0000000000000000; 	// sw
disk[741] <= 32'b010001_11101_01100_0000000100001011; 	// la
disk[742] <= 32'b000000_01100_01011_10011_00000_000000; 	// add
disk[743] <= 32'b001111_11110_01101_1111111111111111; 	// lw
disk[744] <= 32'b010010_10011_01101_0000000000000000; 	// sw
disk[745] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[746] <= 32'b010010_11101_10100_0000000001011111; 	// sw
disk[747] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[748] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[749] <= 32'b010010_11110_00001_0000000000000000; 	// sw
disk[750] <= 32'b010001_11101_00101_0000000100000001; 	// la
disk[751] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[752] <= 32'b000000_00101_00110_01111_00000_000000; 	// add
disk[753] <= 32'b001111_01111_01111_0000000000000000; 	// lw
disk[754] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[755] <= 32'b000000_01111_10001_10000_00000_001101; 	// ne
disk[756] <= 32'b010101_10000_00000_0000001100010111; 	// jf
disk[757] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[758] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[759] <= 32'b100100_00000_00001_0000000000000000; 	// lcdCurr
disk[760] <= 32'b001111_11101_01000_0000000100100001; 	// lw
disk[761] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[762] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[763] <= 32'b001110_11110_10010_0000000000000000; 	// mov
disk[764] <= 32'b000001_10010_10011_0000000000000001; 	// addi
disk[765] <= 32'b010010_11101_10011_0000000010100110; 	// sw
disk[766] <= 32'b010001_11101_01001_0000000000000100; 	// la
disk[767] <= 32'b000000_01001_00110_10100_00000_000000; 	// add
disk[768] <= 32'b001111_11101_01010_0000000000000000; 	// lw
disk[769] <= 32'b010010_10100_01010_0000000000000000; 	// sw
disk[770] <= 32'b010001_11101_01011_0000000000001110; 	// la
disk[771] <= 32'b000000_01011_00110_10101_00000_000000; 	// add
disk[772] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[773] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[774] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[775] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
disk[776] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[777] <= 32'b100000_00000000000000000000000000; 	// exec
disk[778] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[779] <= 32'b010001_11101_00101_0000000000000100; 	// la
disk[780] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[781] <= 32'b000000_00101_00110_10111_00000_000000; 	// add
disk[782] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[783] <= 32'b010010_10111_01111_0000000000000000; 	// sw
disk[784] <= 32'b010001_11101_00111_0000000000001110; 	// la
disk[785] <= 32'b000000_00111_00110_10000_00000_000000; 	// add
disk[786] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[787] <= 32'b010010_10000_10001_0000000000000000; 	// sw
disk[788] <= 32'b001111_11101_01000_0000000100011000; 	// lw
disk[789] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[790] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[791] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[792] <= 32'b000001_11110_11110_0000000000001000; 	// addi
disk[793] <= 32'b010010_11110_00001_1111111111111011; 	// sw
disk[794] <= 32'b001111_11110_00101_1111111111111011; 	// lw
disk[795] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[796] <= 32'b100100_00000_00001_0000000000000000; 	// lcdCurr
disk[797] <= 32'b001111_11101_00110_0000000100100001; 	// lw
disk[798] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[799] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[800] <= 32'b001110_11110_01111_0000000000000000; 	// mov
disk[801] <= 32'b000001_01111_10000_0000000000000001; 	// addi
disk[802] <= 32'b010010_11101_10000_0000000010100110; 	// sw
disk[803] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[804] <= 32'b001111_11101_01000_0000000001011111; 	// lw
disk[805] <= 32'b000000_00111_01000_10001_00000_000000; 	// add
disk[806] <= 32'b001111_11101_01001_0000000000000000; 	// lw
disk[807] <= 32'b010010_10001_01001_0000000000000000; 	// sw
disk[808] <= 32'b010001_11101_01010_0000000001000000; 	// la
disk[809] <= 32'b000000_01010_01000_10010_00000_000000; 	// add
disk[810] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[811] <= 32'b010010_11110_10010_1111111111111101; 	// sw
disk[812] <= 32'b001110_11110_10011_0000000000000000; 	// mov
disk[813] <= 32'b000001_10011_10100_0000000000000001; 	// addi
disk[814] <= 32'b010010_11110_10100_1111111111111110; 	// sw
disk[815] <= 32'b001111_11110_01011_1111111111111101; 	// lw
disk[816] <= 32'b001111_11101_01100_0000000010100000; 	// lw
disk[817] <= 32'b000000_01011_01100_10101_00000_000010; 	// mul
disk[818] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[819] <= 32'b010001_11101_01101_0000000000011000; 	// la
disk[820] <= 32'b000000_01101_01000_10110_00000_000000; 	// add
disk[821] <= 32'b001111_10110_10110_0000000000000000; 	// lw
disk[822] <= 32'b010010_11110_10110_0000000000000000; 	// sw
disk[823] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[824] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[825] <= 32'b000000_00101_01111_10111_00000_010000; 	// gt
disk[826] <= 32'b010101_10111_00000_0000001101001110; 	// jf
disk[827] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[828] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[829] <= 32'b001111_00001_10000_0000000000000000; 	// lw
disk[830] <= 32'b010010_11110_10000_1111111111111100; 	// sw
disk[831] <= 32'b001111_11110_00111_1111111111111100; 	// lw
disk[832] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[833] <= 32'b001111_11110_01000_1111111111111110; 	// lw
disk[834] <= 32'b001110_01000_00010_0000000000000000; 	// mov
disk[835] <= 32'b010010_00010_00001_0000000000000000; 	// sw
disk[836] <= 32'b000001_01000_10001_0000000000000001; 	// addi
disk[837] <= 32'b010010_11110_10001_1111111111111110; 	// sw
disk[838] <= 32'b001111_11110_01000_1111111111111110; 	// lw
disk[839] <= 32'b000001_00110_10010_0000000000000001; 	// addi
disk[840] <= 32'b010010_11110_10010_1111111111111111; 	// sw
disk[841] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[842] <= 32'b000010_00101_10011_0000000000000001; 	// subi
disk[843] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[844] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[845] <= 32'b111100_00000000000000001100110111; 	// j
disk[846] <= 32'b001110_11110_10100_0000000000000000; 	// mov
disk[847] <= 32'b010001_11101_00101_0000000000011000; 	// la
disk[848] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[849] <= 32'b000000_00101_00110_10101_00000_000000; 	// add
disk[850] <= 32'b001111_10101_10101_0000000000000000; 	// lw
disk[851] <= 32'b000000_10100_10101_10110_00000_000000; 	// add
disk[852] <= 32'b001110_10110_00001_0000000000000000; 	// mov
disk[853] <= 32'b001110_00001_11100_0000000000000000; 	// mov
disk[854] <= 32'b000001_00110_10111_0000000000000001; 	// addi
disk[855] <= 32'b001110_10111_00001_0000000000000000; 	// mov
disk[856] <= 32'b010001_11101_00111_0000000000001110; 	// la
disk[857] <= 32'b000000_00111_00110_01111_00000_000000; 	// add
disk[858] <= 32'b001111_01111_01111_0000000000000000; 	// lw
disk[859] <= 32'b001110_01111_00010_0000000000000000; 	// mov
disk[860] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
disk[861] <= 32'b010010_11110_11111_1111111111111010; 	// sw
disk[862] <= 32'b001110_11100_11110_0000000000000000; 	// mov
disk[863] <= 32'b001110_11011_11101_0000000000000000; 	// mov
disk[864] <= 32'b001110_00010_11010_0000000000000000; 	// mov
disk[865] <= 32'b001111_00000_00000_0000011111100000; 	// lw
disk[866] <= 32'b001111_00000_00001_0000011111100001; 	// lw
disk[867] <= 32'b001111_00000_00010_0000011111100010; 	// lw
disk[868] <= 32'b001111_00000_00011_0000011111100011; 	// lw
disk[869] <= 32'b001111_00000_00100_0000011111100100; 	// lw
disk[870] <= 32'b001111_00000_00101_0000011111100101; 	// lw
disk[871] <= 32'b001111_00000_00110_0000011111100110; 	// lw
disk[872] <= 32'b001111_00000_00111_0000011111100111; 	// lw
disk[873] <= 32'b001111_00000_01000_0000011111101000; 	// lw
disk[874] <= 32'b001111_00000_01001_0000011111101001; 	// lw
disk[875] <= 32'b001111_00000_01010_0000011111101010; 	// lw
disk[876] <= 32'b001111_00000_01011_0000011111101011; 	// lw
disk[877] <= 32'b001111_00000_01100_0000011111101100; 	// lw
disk[878] <= 32'b001111_00000_01101_0000011111101101; 	// lw
disk[879] <= 32'b001111_00000_01110_0000011111101110; 	// lw
disk[880] <= 32'b001111_00000_01111_0000011111101111; 	// lw
disk[881] <= 32'b001111_00000_10000_0000011111110000; 	// lw
disk[882] <= 32'b001111_00000_10001_0000011111110001; 	// lw
disk[883] <= 32'b001111_00000_10010_0000011111110010; 	// lw
disk[884] <= 32'b001111_00000_10011_0000011111110011; 	// lw
disk[885] <= 32'b001111_00000_10100_0000011111110100; 	// lw
disk[886] <= 32'b001111_00000_10101_0000011111110101; 	// lw
disk[887] <= 32'b001111_00000_10110_0000011111110110; 	// lw
disk[888] <= 32'b001111_00000_10111_0000011111110111; 	// lw
disk[889] <= 32'b001111_00000_11000_0000011111111000; 	// lw
disk[890] <= 32'b001111_00000_11111_0000011111111001; 	// lw
disk[891] <= 32'b100001_11010_00000_0000000000000000; 	// execAgain
disk[892] <= 32'b001111_11110_11111_1111111111111010; 	// lw
disk[893] <= 32'b010001_11101_00101_0000000000000100; 	// la
disk[894] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[895] <= 32'b000000_00101_00110_10000_00000_000000; 	// add
disk[896] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[897] <= 32'b010010_10000_10001_0000000000000000; 	// sw
disk[898] <= 32'b010001_11101_00111_0000000000001110; 	// la
disk[899] <= 32'b000000_00111_00110_10010_00000_000000; 	// add
disk[900] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[901] <= 32'b010010_10010_10011_0000000000000000; 	// sw
disk[902] <= 32'b001111_11101_01000_0000000100011000; 	// lw
disk[903] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[904] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[905] <= 32'b010000_00000_10100_0000001111100111; 	// li
disk[906] <= 32'b010010_11101_10100_0000000001011110; 	// sw
disk[907] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[908] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[909] <= 32'b010010_11110_00001_1111111111111110; 	// sw
disk[910] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[911] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[912] <= 32'b010010_11110_01111_1111111111111110; 	// sw
disk[913] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[914] <= 32'b010001_11101_00110_0000000011110111; 	// la
disk[915] <= 32'b000000_00110_00101_10000_00000_000000; 	// add
disk[916] <= 32'b001111_10000_10000_0000000000000000; 	// lw
disk[917] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[918] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[919] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[920] <= 32'b010110_00001_10001_0000000000000000; 	// ldk
disk[921] <= 32'b010010_11110_10001_0000000000000000; 	// sw
disk[922] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[923] <= 32'b001101_00101_10010_0000000000011010; 	// srli
disk[924] <= 32'b001111_11101_00110_0000000100010101; 	// lw
disk[925] <= 32'b000000_10010_00110_10011_00000_001101; 	// ne
disk[926] <= 32'b010101_10011_00000_0000001110101011; 	// jf
disk[927] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[928] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[929] <= 32'b001110_00111_00010_0000000000000000; 	// mov
disk[930] <= 32'b010111_00010_00001_0000000000000000; 	// sdk
disk[931] <= 32'b000001_00111_10100_0000000000000001; 	// addi
disk[932] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[933] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[934] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[935] <= 32'b010110_00001_10101_0000000000000000; 	// ldk
disk[936] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[937] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[938] <= 32'b111100_00000000000000001110011010; 	// j
disk[939] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[940] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[941] <= 32'b001110_00101_00010_0000000000000000; 	// mov
disk[942] <= 32'b010111_00010_00001_0000000000000000; 	// sdk
disk[943] <= 32'b010010_11110_11111_1111111111111101; 	// sw
disk[944] <= 32'b111110_00000000000000000011111101; 	// jal
disk[945] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[946] <= 32'b001111_11110_11111_1111111111111101; 	// lw
disk[947] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[948] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[949] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[950] <= 32'b010010_11110_00001_1111111111111110; 	// sw
disk[951] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[952] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[953] <= 32'b010010_11101_01111_0000000001011111; 	// sw
disk[954] <= 32'b010001_11101_00110_0000000000110110; 	// la
disk[955] <= 32'b001111_11101_00111_0000000001011111; 	// lw
disk[956] <= 32'b000000_00110_00111_10000_00000_000000; 	// add
disk[957] <= 32'b001111_10000_10000_0000000000000000; 	// lw
disk[958] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[959] <= 32'b010001_11101_01000_0000000001001010; 	// la
disk[960] <= 32'b000000_01000_00111_10001_00000_000000; 	// add
disk[961] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[962] <= 32'b010010_11110_10001_0000000000000000; 	// sw
disk[963] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[964] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[965] <= 32'b000000_00101_10011_10010_00000_010000; 	// gt
disk[966] <= 32'b010101_10010_00000_0000001111010011; 	// jf
disk[967] <= 32'b010001_11101_00110_0000000001100000; 	// la
disk[968] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[969] <= 32'b000000_00110_00111_10100_00000_000000; 	// add
disk[970] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[971] <= 32'b010010_10100_10101_0000000000000000; 	// sw
disk[972] <= 32'b000001_00111_10110_0000000000000001; 	// addi
disk[973] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[974] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[975] <= 32'b000010_00101_10111_0000000000000001; 	// subi
disk[976] <= 32'b010010_11110_10111_0000000000000000; 	// sw
disk[977] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[978] <= 32'b111100_00000000000000001111000011; 	// j
disk[979] <= 32'b010001_11101_00101_0000000100000001; 	// la
disk[980] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[981] <= 32'b000000_00101_00110_01111_00000_000000; 	// add
disk[982] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[983] <= 32'b010010_01111_10000_0000000000000000; 	// sw
disk[984] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[985] <= 32'b000000_00111_00110_10001_00000_000000; 	// add
disk[986] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[987] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[988] <= 32'b010001_11101_01000_0000000000001110; 	// la
disk[989] <= 32'b000000_01000_00110_10011_00000_000000; 	// add
disk[990] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[991] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[992] <= 32'b010001_11101_01001_0000000000011000; 	// la
disk[993] <= 32'b000000_01001_00110_10101_00000_000000; 	// add
disk[994] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[995] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[996] <= 32'b010001_11101_01010_0000000000100010; 	// la
disk[997] <= 32'b000000_01010_00110_10111_00000_000000; 	// add
disk[998] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[999] <= 32'b010010_10111_01111_0000000000000000; 	// sw
disk[1000] <= 32'b010001_11101_01011_0000000000101100; 	// la
disk[1001] <= 32'b000000_01011_00110_10000_00000_000000; 	// add
disk[1002] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[1003] <= 32'b010010_10000_10001_0000000000000000; 	// sw
disk[1004] <= 32'b010001_11101_01100_0000000001000000; 	// la
disk[1005] <= 32'b000000_01100_00110_10010_00000_000000; 	// add
disk[1006] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[1007] <= 32'b010010_10010_10011_0000000000000000; 	// sw
disk[1008] <= 32'b010001_11101_01101_0000000001001010; 	// la
disk[1009] <= 32'b000000_01101_00110_10100_00000_000000; 	// add
disk[1010] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[1011] <= 32'b010010_10100_10101_0000000000000000; 	// sw
disk[1012] <= 32'b010001_11101_01110_0000000001010100; 	// la
disk[1013] <= 32'b000000_01110_00110_10110_00000_000000; 	// add
disk[1014] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[1015] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[1016] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[1017] <= 32'b010010_11101_01111_0000000001011111; 	// sw
disk[1018] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[1019] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[1020] <= 32'b000001_11110_11110_0000000000000111; 	// addi
disk[1021] <= 32'b010010_11110_00001_1111111111111100; 	// sw
disk[1022] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[1023] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[1024] <= 32'b010010_11101_01111_0000000001011111; 	// sw
disk[1025] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[1026] <= 32'b010010_11101_00110_0000000001011110; 	// sw
disk[1027] <= 32'b010001_11101_00111_0000000001000000; 	// la
disk[1028] <= 32'b000000_00111_00110_10000_00000_000000; 	// add
disk[1029] <= 32'b001111_10000_10000_0000000000000000; 	// lw
disk[1030] <= 32'b000001_10000_10001_0000000000000001; 	// addi
disk[1031] <= 32'b010010_11110_10001_1111111111111110; 	// sw
disk[1032] <= 32'b001111_11110_01000_1111111111111110; 	// lw
disk[1033] <= 32'b001111_11101_01001_0000000010100000; 	// lw
disk[1034] <= 32'b000000_01000_01001_10010_00000_000010; 	// mul
disk[1035] <= 32'b010010_11110_10010_1111111111111111; 	// sw
disk[1036] <= 32'b001111_11101_01010_0000000010100001; 	// lw
disk[1037] <= 32'b000010_01010_10011_0000000000000001; 	// subi
disk[1038] <= 32'b000000_01001_10011_10100_00000_000010; 	// mul
disk[1039] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[1040] <= 32'b001111_11101_00101_0000000010100000; 	// lw
disk[1041] <= 32'b001111_11101_00110_0000000010100001; 	// lw
disk[1042] <= 32'b000000_00101_00110_10101_00000_000010; 	// mul
disk[1043] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[1044] <= 32'b000000_00111_10101_10110_00000_001110; 	// lt
disk[1045] <= 32'b010101_10110_00000_0000010000100101; 	// jf
disk[1046] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[1047] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[1048] <= 32'b001111_00001_10111_0000000000000000; 	// lw
disk[1049] <= 32'b010010_11110_10111_1111111111111101; 	// sw
disk[1050] <= 32'b001111_11110_01001_1111111111111101; 	// lw
disk[1051] <= 32'b001110_01001_00001_0000000000000000; 	// mov
disk[1052] <= 32'b001110_00111_00010_0000000000000000; 	// mov
disk[1053] <= 32'b010010_00010_00001_0000000000000000; 	// sw
disk[1054] <= 32'b000001_01000_01111_0000000000000001; 	// addi
disk[1055] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[1056] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[1057] <= 32'b000001_00111_10000_0000000000000001; 	// addi
disk[1058] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[1059] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[1060] <= 32'b111100_00000000000000010000010000; 	// j
disk[1061] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[1062] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1063] <= 32'b010010_11110_11111_1111111111111011; 	// sw
disk[1064] <= 32'b111110_00000000000000001100011000; 	// jal
disk[1065] <= 32'b000010_11110_11110_0000000000001000; 	// subi
disk[1066] <= 32'b001111_11110_11111_1111111111111011; 	// lw
disk[1067] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1068] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[1069] <= 32'b010000_00000_11110_0000000100101001; 	// li
disk[1070] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[1071] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[1072] <= 32'b010010_11110_00001_0000000000000000; 	// sw
disk[1073] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1074] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[1075] <= 32'b010010_11101_01111_0000000001011111; 	// sw
disk[1076] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[1077] <= 32'b010010_11101_00110_0000000001011110; 	// sw
disk[1078] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1079] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[1080] <= 32'b111110_00000000000000001011101100; 	// jal
disk[1081] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1082] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[1083] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1084] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[1085] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[1086] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[1087] <= 32'b111110_00000000000000001001100001; 	// jal
disk[1088] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1089] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[1090] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1091] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[1092] <= 32'b111110_00000000000000001001001010; 	// jal
disk[1093] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1094] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[1095] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1096] <= 32'b001111_11101_00110_0000000000000011; 	// lw
disk[1097] <= 32'b000000_00101_00110_01111_00000_001101; 	// ne
disk[1098] <= 32'b010101_01111_00000_0000010001011010; 	// jf
disk[1099] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[1100] <= 32'b111110_00000000000000001001001010; 	// jal
disk[1101] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1102] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[1103] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1104] <= 32'b010010_11101_00101_0000000001011111; 	// sw
disk[1105] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[1106] <= 32'b000001_00110_10000_0000000000000001; 	// addi
disk[1107] <= 32'b001110_10000_00001_0000000000000000; 	// mov
disk[1108] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[1109] <= 32'b111110_00000000000000001011101100; 	// jal
disk[1110] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1111] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[1112] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1113] <= 32'b111100_00000000000000010001000011; 	// j
disk[1114] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[1115] <= 32'b001110_11110_11100_0000000000000000; 	// mov
disk[1116] <= 32'b001110_11101_11011_0000000000000000; 	// mov
disk[1117] <= 32'b010000_00000_00000_0000000000000000; 	// li
disk[1118] <= 32'b010000_00000_11110_0000000000000000; 	// li
disk[1119] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[1120] <= 32'b000001_11110_11110_0000000100101100; 	// addi
disk[1121] <= 32'b010010_00000_00000_0000011111100000; 	// sw
disk[1122] <= 32'b010010_00000_00001_0000011111100001; 	// sw
disk[1123] <= 32'b010010_00000_00010_0000011111100010; 	// sw
disk[1124] <= 32'b010010_00000_00011_0000011111100011; 	// sw
disk[1125] <= 32'b010010_00000_00100_0000011111100100; 	// sw
disk[1126] <= 32'b010010_00000_00101_0000011111100101; 	// sw
disk[1127] <= 32'b010010_00000_00110_0000011111100110; 	// sw
disk[1128] <= 32'b010010_00000_00111_0000011111100111; 	// sw
disk[1129] <= 32'b010010_00000_01000_0000011111101000; 	// sw
disk[1130] <= 32'b010010_00000_01001_0000011111101001; 	// sw
disk[1131] <= 32'b010010_00000_01010_0000011111101010; 	// sw
disk[1132] <= 32'b010010_00000_01011_0000011111101011; 	// sw
disk[1133] <= 32'b010010_00000_01100_0000011111101100; 	// sw
disk[1134] <= 32'b010010_00000_01101_0000011111101101; 	// sw
disk[1135] <= 32'b010010_00000_01110_0000011111101110; 	// sw
disk[1136] <= 32'b010010_00000_01111_0000011111101111; 	// sw
disk[1137] <= 32'b010010_00000_10000_0000011111110000; 	// sw
disk[1138] <= 32'b010010_00000_10001_0000011111110001; 	// sw
disk[1139] <= 32'b010010_00000_10010_0000011111110010; 	// sw
disk[1140] <= 32'b010010_00000_10011_0000011111110011; 	// sw
disk[1141] <= 32'b010010_00000_10100_0000011111110100; 	// sw
disk[1142] <= 32'b010010_00000_10101_0000011111110101; 	// sw
disk[1143] <= 32'b010010_00000_10110_0000011111110110; 	// sw
disk[1144] <= 32'b010010_00000_10111_0000011111110111; 	// sw
disk[1145] <= 32'b010010_00000_11000_0000011111111000; 	// sw
disk[1146] <= 32'b010010_00000_11111_0000011111111001; 	// sw
disk[1147] <= 32'b001111_11110_00101_1111111111111011; 	// lw
disk[1148] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[1149] <= 32'b000000_00101_10000_01111_00000_001100; 	// eq
disk[1150] <= 32'b010101_01111_00000_0000010010001000; 	// jf
disk[1151] <= 32'b111110_00000000000000000100111001; 	// jal
disk[1152] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[1153] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1154] <= 32'b001111_11101_00110_0000000100011000; 	// lw
disk[1155] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1156] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[1157] <= 32'b010000_00000_10001_0000000000000001; 	// li
disk[1158] <= 32'b010010_11110_10001_1111111111111011; 	// sw
disk[1159] <= 32'b100110_00000_00000_0000000000000000; 	// cic
disk[1160] <= 32'b100101_00000_10010_0000000000000000; 	// gic
disk[1161] <= 32'b010010_11110_10010_1111111111111010; 	// sw
disk[1162] <= 32'b001111_11110_00101_1111111111111010; 	// lw
disk[1163] <= 32'b010000_00000_10100_0000000000000001; 	// li
disk[1164] <= 32'b000000_00101_10100_10011_00000_001100; 	// eq
disk[1165] <= 32'b010101_10011_00000_0000010100001100; 	// jf
disk[1166] <= 32'b001110_11100_10101_0000000000000000; 	// mov
disk[1167] <= 32'b010010_11101_10101_0000000010100111; 	// sw
disk[1168] <= 32'b001111_11101_00110_0000000010100111; 	// lw
disk[1169] <= 32'b001111_11101_00111_0000000010100110; 	// lw
disk[1170] <= 32'b000000_00110_00111_10110_00000_000001; 	// sub
disk[1171] <= 32'b000001_10110_10111_0000000000000001; 	// addi
disk[1172] <= 32'b010010_11110_10111_0000000000000000; 	// sw
disk[1173] <= 32'b010001_11101_01000_0000000000011000; 	// la
disk[1174] <= 32'b001111_11101_01001_0000000001011111; 	// lw
disk[1175] <= 32'b000000_01000_01001_01111_00000_000000; 	// add
disk[1176] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[1177] <= 32'b010010_01111_01010_0000000000000000; 	// sw
disk[1178] <= 32'b010001_11101_01011_0000000000000100; 	// la
disk[1179] <= 32'b000000_01011_01001_10000_00000_000000; 	// add
disk[1180] <= 32'b001111_11101_01100_0000000000000010; 	// lw
disk[1181] <= 32'b010010_10000_01100_0000000000000000; 	// sw
disk[1182] <= 32'b100111_00000_10001_0000000000000000; 	// gip
disk[1183] <= 32'b000001_10001_10010_0000000000000001; 	// addi
disk[1184] <= 32'b010001_11101_01101_0000000000001110; 	// la
disk[1185] <= 32'b000000_01101_01001_10011_00000_000000; 	// add
disk[1186] <= 32'b010010_10011_10010_0000000000000000; 	// sw
disk[1187] <= 32'b010001_11101_01110_0000000001000000; 	// la
disk[1188] <= 32'b000000_01110_01001_10100_00000_000000; 	// add
disk[1189] <= 32'b001111_10100_10100_0000000000000000; 	// lw
disk[1190] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[1191] <= 32'b000000_10100_10110_10101_00000_001100; 	// eq
disk[1192] <= 32'b010101_10101_00000_0000010010110011; 	// jf
disk[1193] <= 32'b111110_00000000000000000110010100; 	// jal
disk[1194] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[1195] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1196] <= 32'b010010_11110_00101_1111111111111100; 	// sw
disk[1197] <= 32'b010001_11101_00110_0000000001000000; 	// la
disk[1198] <= 32'b001111_11101_00111_0000000001011111; 	// lw
disk[1199] <= 32'b000000_00110_00111_10111_00000_000000; 	// add
disk[1200] <= 32'b001111_11110_01000_1111111111111100; 	// lw
disk[1201] <= 32'b010010_10111_01000_0000000000000000; 	// sw
disk[1202] <= 32'b111100_00000000000000010010111000; 	// j
disk[1203] <= 32'b010001_11101_00101_0000000001000000; 	// la
disk[1204] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[1205] <= 32'b000000_00101_00110_01111_00000_000000; 	// add
disk[1206] <= 32'b001111_01111_01111_0000000000000000; 	// lw
disk[1207] <= 32'b010010_11110_01111_1111111111111100; 	// sw
disk[1208] <= 32'b001111_11101_00101_0000000010100110; 	// lw
disk[1209] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[1210] <= 32'b001111_11110_00110_1111111111111100; 	// lw
disk[1211] <= 32'b001111_11101_00111_0000000010100000; 	// lw
disk[1212] <= 32'b000000_00110_00111_10000_00000_000010; 	// mul
disk[1213] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[1214] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1215] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[1216] <= 32'b000000_00101_10010_10001_00000_010000; 	// gt
disk[1217] <= 32'b010101_10001_00000_0000010011010101; 	// jf
disk[1218] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[1219] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1220] <= 32'b001111_00001_10011_0000000000000000; 	// lw
disk[1221] <= 32'b010010_11110_10011_1111111111111101; 	// sw
disk[1222] <= 32'b001111_11110_00111_1111111111111101; 	// lw
disk[1223] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1224] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[1225] <= 32'b001110_01000_00010_0000000000000000; 	// mov
disk[1226] <= 32'b010010_00010_00001_0000000000000000; 	// sw
disk[1227] <= 32'b000001_00110_10100_0000000000000001; 	// addi
disk[1228] <= 32'b010010_11110_10100_1111111111111110; 	// sw
disk[1229] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[1230] <= 32'b000001_01000_10101_0000000000000001; 	// addi
disk[1231] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[1232] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[1233] <= 32'b000010_00101_10110_0000000000000001; 	// subi
disk[1234] <= 32'b010010_11110_10110_0000000000000000; 	// sw
disk[1235] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1236] <= 32'b111100_00000000000000010010111110; 	// j
disk[1237] <= 32'b001111_11101_00101_0000000001011111; 	// lw
disk[1238] <= 32'b001111_11101_00110_0000000001011110; 	// lw
disk[1239] <= 32'b000000_00101_00110_10111_00000_001100; 	// eq
disk[1240] <= 32'b010101_10111_00000_0000010011100000; 	// jf
disk[1241] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1242] <= 32'b111110_00000000000000001100011000; 	// jal
disk[1243] <= 32'b000010_11110_11110_0000000000001000; 	// subi
disk[1244] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1245] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[1246] <= 32'b010000_00000_11110_0000000100101100; 	// li
disk[1247] <= 32'b111100_00000000000000010100000101; 	// j
disk[1248] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[1249] <= 32'b000001_00101_01111_0000000000000001; 	// addi
disk[1250] <= 32'b010010_11110_01111_1111111111111100; 	// sw
disk[1251] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[1252] <= 32'b001111_11101_00110_0000000010100001; 	// lw
disk[1253] <= 32'b000010_00110_10000_0000000000000001; 	// subi
disk[1254] <= 32'b001111_11101_00111_0000000010100000; 	// lw
disk[1255] <= 32'b000000_00111_10000_10001_00000_000010; 	// mul
disk[1256] <= 32'b010010_11110_10001_1111111111111110; 	// sw
disk[1257] <= 32'b000000_00101_00111_10010_00000_000010; 	// mul
disk[1258] <= 32'b010010_11110_10010_1111111111111111; 	// sw
disk[1259] <= 32'b001111_11101_00101_0000000010100000; 	// lw
disk[1260] <= 32'b001111_11101_00110_0000000010100001; 	// lw
disk[1261] <= 32'b000000_00101_00110_10011_00000_000010; 	// mul
disk[1262] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[1263] <= 32'b000000_00111_10011_10100_00000_001110; 	// lt
disk[1264] <= 32'b010101_10100_00000_0000010100000000; 	// jf
disk[1265] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1266] <= 32'b001111_00001_10101_0000000000000000; 	// lw
disk[1267] <= 32'b010010_11110_10101_1111111111111101; 	// sw
disk[1268] <= 32'b001111_11110_01000_1111111111111101; 	// lw
disk[1269] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[1270] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[1271] <= 32'b001110_01001_00010_0000000000000000; 	// mov
disk[1272] <= 32'b010010_00010_00001_0000000000000000; 	// sw
disk[1273] <= 32'b000001_00111_10110_0000000000000001; 	// addi
disk[1274] <= 32'b010010_11110_10110_1111111111111110; 	// sw
disk[1275] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[1276] <= 32'b000001_01001_10111_0000000000000001; 	// addi
disk[1277] <= 32'b010010_11110_10111_1111111111111111; 	// sw
disk[1278] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[1279] <= 32'b111100_00000000000000010011101011; 	// j
disk[1280] <= 32'b010001_11101_00101_0000000000000100; 	// la
disk[1281] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[1282] <= 32'b000000_00101_00110_01111_00000_000000; 	// add
disk[1283] <= 32'b001111_11101_00111_0000000000000010; 	// lw
disk[1284] <= 32'b010010_01111_00111_0000000000000000; 	// sw
disk[1285] <= 32'b001111_11101_00101_0000000100011000; 	// lw
disk[1286] <= 32'b010010_11101_00101_0000000100100010; 	// sw
disk[1287] <= 32'b001111_11101_00110_0000000100100010; 	// lw
disk[1288] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1289] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[1290] <= 32'b100110_00000_00000_0000000000000000; 	// cic
disk[1291] <= 32'b111100_00000000000000010110000001; 	// j
disk[1292] <= 32'b001111_11110_00101_1111111111111010; 	// lw
disk[1293] <= 32'b010000_00000_10001_0000000000000010; 	// li
disk[1294] <= 32'b000000_00101_10001_10000_00000_001100; 	// eq
disk[1295] <= 32'b010101_10000_00000_0000010110000001; 	// jf
disk[1296] <= 32'b001110_11100_10010_0000000000000000; 	// mov
disk[1297] <= 32'b010010_11101_10010_0000000010100111; 	// sw
disk[1298] <= 32'b001111_11101_00110_0000000010100111; 	// lw
disk[1299] <= 32'b001111_11101_00111_0000000010100110; 	// lw
disk[1300] <= 32'b000000_00110_00111_10011_00000_000001; 	// sub
disk[1301] <= 32'b000001_10011_10100_0000000000000001; 	// addi
disk[1302] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[1303] <= 32'b010001_11101_01000_0000000000011000; 	// la
disk[1304] <= 32'b001111_11101_01001_0000000001011111; 	// lw
disk[1305] <= 32'b000000_01000_01001_10101_00000_000000; 	// add
disk[1306] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[1307] <= 32'b010010_10101_01010_0000000000000000; 	// sw
disk[1308] <= 32'b010001_11101_01011_0000000000000100; 	// la
disk[1309] <= 32'b000000_01011_01001_10110_00000_000000; 	// add
disk[1310] <= 32'b001111_11101_01100_0000000000000010; 	// lw
disk[1311] <= 32'b010010_10110_01100_0000000000000000; 	// sw
disk[1312] <= 32'b100111_00000_10111_0000000000000000; 	// gip
disk[1313] <= 32'b010001_11101_01101_0000000000001110; 	// la
disk[1314] <= 32'b000000_01101_01001_01111_00000_000000; 	// add
disk[1315] <= 32'b010010_01111_10111_0000000000000000; 	// sw
disk[1316] <= 32'b010001_11101_01110_0000000001000000; 	// la
disk[1317] <= 32'b000000_01110_01001_10000_00000_000000; 	// add
disk[1318] <= 32'b001111_10000_10000_0000000000000000; 	// lw
disk[1319] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[1320] <= 32'b000000_10000_10010_10001_00000_001100; 	// eq
disk[1321] <= 32'b010101_10001_00000_0000010100110100; 	// jf
disk[1322] <= 32'b111110_00000000000000000110010100; 	// jal
disk[1323] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[1324] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1325] <= 32'b010010_11110_00101_1111111111111100; 	// sw
disk[1326] <= 32'b010001_11101_00110_0000000001000000; 	// la
disk[1327] <= 32'b001111_11101_00111_0000000001011111; 	// lw
disk[1328] <= 32'b000000_00110_00111_10011_00000_000000; 	// add
disk[1329] <= 32'b001111_11110_01000_1111111111111100; 	// lw
disk[1330] <= 32'b010010_10011_01000_0000000000000000; 	// sw
disk[1331] <= 32'b111100_00000000000000010100111001; 	// j
disk[1332] <= 32'b010001_11101_00101_0000000001000000; 	// la
disk[1333] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[1334] <= 32'b000000_00101_00110_10100_00000_000000; 	// add
disk[1335] <= 32'b001111_10100_10100_0000000000000000; 	// lw
disk[1336] <= 32'b010010_11110_10100_1111111111111100; 	// sw
disk[1337] <= 32'b001111_11101_00101_0000000010100110; 	// lw
disk[1338] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[1339] <= 32'b001111_11110_00110_1111111111111100; 	// lw
disk[1340] <= 32'b001111_11101_00111_0000000010100000; 	// lw
disk[1341] <= 32'b000000_00110_00111_10101_00000_000010; 	// mul
disk[1342] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[1343] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1344] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[1345] <= 32'b000000_00101_10111_10110_00000_010000; 	// gt
disk[1346] <= 32'b010101_10110_00000_0000010101010110; 	// jf
disk[1347] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[1348] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1349] <= 32'b001111_00001_01111_0000000000000000; 	// lw
disk[1350] <= 32'b010010_11110_01111_1111111111111101; 	// sw
disk[1351] <= 32'b001111_11110_00111_1111111111111101; 	// lw
disk[1352] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1353] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[1354] <= 32'b001110_01000_00010_0000000000000000; 	// mov
disk[1355] <= 32'b010010_00010_00001_0000000000000000; 	// sw
disk[1356] <= 32'b000001_00110_10000_0000000000000001; 	// addi
disk[1357] <= 32'b010010_11110_10000_1111111111111110; 	// sw
disk[1358] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[1359] <= 32'b000001_01000_10001_0000000000000001; 	// addi
disk[1360] <= 32'b010010_11110_10001_1111111111111111; 	// sw
disk[1361] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[1362] <= 32'b000010_00101_10010_0000000000000001; 	// subi
disk[1363] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[1364] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1365] <= 32'b111100_00000000000000010100111111; 	// j
disk[1366] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[1367] <= 32'b000001_00101_10011_0000000000000001; 	// addi
disk[1368] <= 32'b010010_11110_10011_1111111111111100; 	// sw
disk[1369] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[1370] <= 32'b001111_11101_00110_0000000010100001; 	// lw
disk[1371] <= 32'b000010_00110_10100_0000000000000001; 	// subi
disk[1372] <= 32'b001111_11101_00111_0000000010100000; 	// lw
disk[1373] <= 32'b000000_00111_10100_10101_00000_000010; 	// mul
disk[1374] <= 32'b010010_11110_10101_1111111111111110; 	// sw
disk[1375] <= 32'b000000_00101_00111_10110_00000_000010; 	// mul
disk[1376] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[1377] <= 32'b001111_11101_00101_0000000010100000; 	// lw
disk[1378] <= 32'b001111_11101_00110_0000000010100001; 	// lw
disk[1379] <= 32'b000000_00101_00110_10111_00000_000010; 	// mul
disk[1380] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[1381] <= 32'b000000_00111_10111_01111_00000_001110; 	// lt
disk[1382] <= 32'b010101_01111_00000_0000010101110110; 	// jf
disk[1383] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1384] <= 32'b001111_00001_10000_0000000000000000; 	// lw
disk[1385] <= 32'b010010_11110_10000_1111111111111101; 	// sw
disk[1386] <= 32'b001111_11110_01000_1111111111111101; 	// lw
disk[1387] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[1388] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[1389] <= 32'b001110_01001_00010_0000000000000000; 	// mov
disk[1390] <= 32'b010010_00010_00001_0000000000000000; 	// sw
disk[1391] <= 32'b000001_00111_10001_0000000000000001; 	// addi
disk[1392] <= 32'b010010_11110_10001_1111111111111110; 	// sw
disk[1393] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[1394] <= 32'b000001_01001_10010_0000000000000001; 	// addi
disk[1395] <= 32'b010010_11110_10010_1111111111111111; 	// sw
disk[1396] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[1397] <= 32'b111100_00000000000000010101100001; 	// j
disk[1398] <= 32'b010001_11101_00101_0000000000000100; 	// la
disk[1399] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[1400] <= 32'b000000_00101_00110_10011_00000_000000; 	// add
disk[1401] <= 32'b001111_11101_00111_0000000000000010; 	// lw
disk[1402] <= 32'b010010_10011_00111_0000000000000000; 	// sw
disk[1403] <= 32'b001111_11101_01000_0000000100011000; 	// lw
disk[1404] <= 32'b010010_11101_01000_0000000100100010; 	// sw
disk[1405] <= 32'b001111_11101_01001_0000000100100010; 	// lw
disk[1406] <= 32'b001110_01001_00001_0000000000000000; 	// mov
disk[1407] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[1408] <= 32'b100110_00000_00000_0000000000000000; 	// cic
disk[1409] <= 32'b010000_00000_10100_0000000000000001; 	// li
disk[1410] <= 32'b010101_10100_00000_0000011001111010; 	// jf
disk[1411] <= 32'b010011_00000_10101_0000000000000000; 	// in
disk[1412] <= 32'b010010_11110_10101_1111111111111001; 	// sw
disk[1413] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1414] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1415] <= 32'b010000_00000_00010_0000000000000000; 	// li
disk[1416] <= 32'b010100_00000_00001_0000000000000000; 	// out
disk[1417] <= 32'b001111_11101_00110_0000000100100010; 	// lw
disk[1418] <= 32'b001111_11101_00111_0000000100011000; 	// lw
disk[1419] <= 32'b000000_00110_00111_10110_00000_001100; 	// eq
disk[1420] <= 32'b010101_10110_00000_0000010110110001; 	// jf
disk[1421] <= 32'b010000_00000_01111_0000000000000001; 	// li
disk[1422] <= 32'b000000_00101_01111_10111_00000_001100; 	// eq
disk[1423] <= 32'b010101_10111_00000_0000010110010100; 	// jf
disk[1424] <= 32'b001111_11101_01000_0000000100011001; 	// lw
disk[1425] <= 32'b010010_11110_01000_1111111111111001; 	// sw
disk[1426] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1427] <= 32'b111100_00000000000000010110110000; 	// j
disk[1428] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1429] <= 32'b010000_00000_10001_0000000000000010; 	// li
disk[1430] <= 32'b000000_00101_10001_10000_00000_001100; 	// eq
disk[1431] <= 32'b010101_10000_00000_0000010110011100; 	// jf
disk[1432] <= 32'b001111_11101_00110_0000000100011011; 	// lw
disk[1433] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1434] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1435] <= 32'b111100_00000000000000010110110000; 	// j
disk[1436] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1437] <= 32'b010000_00000_10011_0000000000000011; 	// li
disk[1438] <= 32'b000000_00101_10011_10010_00000_001100; 	// eq
disk[1439] <= 32'b010101_10010_00000_0000010110100100; 	// jf
disk[1440] <= 32'b001111_11101_00110_0000000100011110; 	// lw
disk[1441] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1442] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1443] <= 32'b111100_00000000000000010110110000; 	// j
disk[1444] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1445] <= 32'b010000_00000_10101_0000000000000100; 	// li
disk[1446] <= 32'b000000_00101_10101_10100_00000_001100; 	// eq
disk[1447] <= 32'b010101_10100_00000_0000010110101110; 	// jf
disk[1448] <= 32'b111110_00000000000000000000110011; 	// jal
disk[1449] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[1450] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1451] <= 32'b001111_11101_00110_0000000100011000; 	// lw
disk[1452] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1453] <= 32'b111100_00000000000000010110110000; 	// j
disk[1454] <= 32'b001111_11101_00101_0000000100011000; 	// lw
disk[1455] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1456] <= 32'b111100_00000000000000011001110100; 	// j
disk[1457] <= 32'b001111_11101_00101_0000000100100010; 	// lw
disk[1458] <= 32'b001111_11101_00110_0000000100011001; 	// lw
disk[1459] <= 32'b000000_00101_00110_10110_00000_001100; 	// eq
disk[1460] <= 32'b010101_10110_00000_0000010111010101; 	// jf
disk[1461] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1462] <= 32'b010000_00000_01111_0000000000000001; 	// li
disk[1463] <= 32'b000000_00111_01111_10111_00000_001100; 	// eq
disk[1464] <= 32'b010101_10111_00000_0000010110111101; 	// jf
disk[1465] <= 32'b001111_11101_01000_0000000100011000; 	// lw
disk[1466] <= 32'b010010_11110_01000_1111111111111001; 	// sw
disk[1467] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1468] <= 32'b111100_00000000000000010111010100; 	// j
disk[1469] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1470] <= 32'b010000_00000_10001_0000000000000010; 	// li
disk[1471] <= 32'b000000_00101_10001_10000_00000_001100; 	// eq
disk[1472] <= 32'b010101_10000_00000_0000010111000101; 	// jf
disk[1473] <= 32'b001111_11101_00110_0000000100011000; 	// lw
disk[1474] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1475] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1476] <= 32'b111100_00000000000000010111010100; 	// j
disk[1477] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1478] <= 32'b010000_00000_10011_0000000000000011; 	// li
disk[1479] <= 32'b000000_00101_10011_10010_00000_001100; 	// eq
disk[1480] <= 32'b010101_10010_00000_0000010111010010; 	// jf
disk[1481] <= 32'b001111_11101_00110_0000000100011010; 	// lw
disk[1482] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1483] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1484] <= 32'b111110_00000000000000000111110001; 	// jal
disk[1485] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1486] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1487] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1488] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[1489] <= 32'b111100_00000000000000010111010100; 	// j
disk[1490] <= 32'b001111_11101_00101_0000000100011000; 	// lw
disk[1491] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1492] <= 32'b111100_00000000000000011001110100; 	// j
disk[1493] <= 32'b001111_11101_00101_0000000100100010; 	// lw
disk[1494] <= 32'b001111_11101_00110_0000000100011010; 	// lw
disk[1495] <= 32'b000000_00101_00110_10100_00000_001100; 	// eq
disk[1496] <= 32'b010101_10100_00000_0000010111100100; 	// jf
disk[1497] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1498] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[1499] <= 32'b000000_00111_10110_10101_00000_010000; 	// gt
disk[1500] <= 32'b010101_10101_00000_0000010111100001; 	// jf
disk[1501] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1502] <= 32'b111110_00000000000000001110001100; 	// jal
disk[1503] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[1504] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1505] <= 32'b001111_11101_00101_0000000100011000; 	// lw
disk[1506] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1507] <= 32'b111100_00000000000000011001110100; 	// j
disk[1508] <= 32'b001111_11101_00101_0000000100100010; 	// lw
disk[1509] <= 32'b001111_11101_00110_0000000100011011; 	// lw
disk[1510] <= 32'b000000_00101_00110_10111_00000_001100; 	// eq
disk[1511] <= 32'b010101_10111_00000_0000011000010010; 	// jf
disk[1512] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1513] <= 32'b010000_00000_10000_0000000000000001; 	// li
disk[1514] <= 32'b000000_00111_10000_01111_00000_001100; 	// eq
disk[1515] <= 32'b010101_01111_00000_0000010111110101; 	// jf
disk[1516] <= 32'b001111_11101_01000_0000000100011100; 	// lw
disk[1517] <= 32'b010010_11110_01000_1111111111111001; 	// sw
disk[1518] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1519] <= 32'b111110_00000000000000000111110001; 	// jal
disk[1520] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1521] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1522] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1523] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[1524] <= 32'b111100_00000000000000011000010001; 	// j
disk[1525] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1526] <= 32'b010000_00000_10010_0000000000000011; 	// li
disk[1527] <= 32'b000000_00101_10010_10001_00000_001100; 	// eq
disk[1528] <= 32'b010101_10001_00000_0000011000000010; 	// jf
disk[1529] <= 32'b001111_11101_00110_0000000100011101; 	// lw
disk[1530] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1531] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1532] <= 32'b111110_00000000000000000111010000; 	// jal
disk[1533] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1534] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1535] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1536] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[1537] <= 32'b111100_00000000000000011000010001; 	// j
disk[1538] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1539] <= 32'b010000_00000_10100_0000000000000011; 	// li
disk[1540] <= 32'b000000_00101_10100_10011_00000_010000; 	// gt
disk[1541] <= 32'b010101_10011_00000_0000011000001010; 	// jf
disk[1542] <= 32'b001111_11101_00110_0000000100011000; 	// lw
disk[1543] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1544] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1545] <= 32'b111100_00000000000000011000010001; 	// j
disk[1546] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1547] <= 32'b010000_00000_10110_0000000000000001; 	// li
disk[1548] <= 32'b000000_00101_10110_10101_00000_001110; 	// lt
disk[1549] <= 32'b010101_10101_00000_0000011000010001; 	// jf
disk[1550] <= 32'b001111_11101_00110_0000000100011000; 	// lw
disk[1551] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1552] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1553] <= 32'b111100_00000000000000011001110100; 	// j
disk[1554] <= 32'b001111_11101_00101_0000000100100010; 	// lw
disk[1555] <= 32'b001111_11101_00110_0000000100011100; 	// lw
disk[1556] <= 32'b000000_00101_00110_10111_00000_001100; 	// eq
disk[1557] <= 32'b010101_10111_00000_0000011000100001; 	// jf
disk[1558] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1559] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[1560] <= 32'b000000_00111_10000_01111_00000_010000; 	// gt
disk[1561] <= 32'b010101_01111_00000_0000011000011110; 	// jf
disk[1562] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1563] <= 32'b111110_00000000000000001010010011; 	// jal
disk[1564] <= 32'b000010_11110_11110_0000000000001010; 	// subi
disk[1565] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1566] <= 32'b001111_11101_00101_0000000100011000; 	// lw
disk[1567] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1568] <= 32'b111100_00000000000000011001110100; 	// j
disk[1569] <= 32'b001111_11101_00101_0000000100100010; 	// lw
disk[1570] <= 32'b001111_11101_00110_0000000100011101; 	// lw
disk[1571] <= 32'b000000_00101_00110_10001_00000_001100; 	// eq
disk[1572] <= 32'b010101_10001_00000_0000011000110000; 	// jf
disk[1573] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1574] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[1575] <= 32'b000000_00111_10011_10010_00000_010000; 	// gt
disk[1576] <= 32'b010101_10010_00000_0000011000101101; 	// jf
disk[1577] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1578] <= 32'b111110_00000000000000001110110101; 	// jal
disk[1579] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[1580] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1581] <= 32'b001111_11101_00101_0000000100011000; 	// lw
disk[1582] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1583] <= 32'b111100_00000000000000011001110100; 	// j
disk[1584] <= 32'b001111_11101_00101_0000000100100010; 	// lw
disk[1585] <= 32'b001111_11101_00110_0000000100011110; 	// lw
disk[1586] <= 32'b000000_00101_00110_10100_00000_001100; 	// eq
disk[1587] <= 32'b010101_10100_00000_0000011001011001; 	// jf
disk[1588] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1589] <= 32'b010000_00000_10110_0000000000000001; 	// li
disk[1590] <= 32'b000000_00111_10110_10101_00000_001100; 	// eq
disk[1591] <= 32'b010101_10101_00000_0000011000111110; 	// jf
disk[1592] <= 32'b111110_00000000000000010000111101; 	// jal
disk[1593] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[1594] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1595] <= 32'b001111_11101_00110_0000000100011000; 	// lw
disk[1596] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1597] <= 32'b111100_00000000000000011001011000; 	// j
disk[1598] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1599] <= 32'b010000_00000_01111_0000000000000010; 	// li
disk[1600] <= 32'b000000_00101_01111_10111_00000_001100; 	// eq
disk[1601] <= 32'b010101_10111_00000_0000011001001010; 	// jf
disk[1602] <= 32'b111110_00000000000000000111010000; 	// jal
disk[1603] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1604] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1605] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1606] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[1607] <= 32'b001111_11101_00110_0000000100011111; 	// lw
disk[1608] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1609] <= 32'b111100_00000000000000011001011000; 	// j
disk[1610] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1611] <= 32'b010000_00000_10001_0000000000000011; 	// li
disk[1612] <= 32'b000000_00101_10001_10000_00000_001100; 	// eq
disk[1613] <= 32'b010101_10000_00000_0000011001010110; 	// jf
disk[1614] <= 32'b111110_00000000000000001000010010; 	// jal
disk[1615] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1616] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1617] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1618] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[1619] <= 32'b001111_11101_00110_0000000100100000; 	// lw
disk[1620] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1621] <= 32'b111100_00000000000000011001011000; 	// j
disk[1622] <= 32'b001111_11101_00101_0000000100011000; 	// lw
disk[1623] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1624] <= 32'b111100_00000000000000011001110100; 	// j
disk[1625] <= 32'b001111_11101_00101_0000000100100010; 	// lw
disk[1626] <= 32'b001111_11101_00110_0000000100011111; 	// lw
disk[1627] <= 32'b000000_00101_00110_10010_00000_001100; 	// eq
disk[1628] <= 32'b010101_10010_00000_0000011001101000; 	// jf
disk[1629] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1630] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[1631] <= 32'b000000_00111_10100_10011_00000_010000; 	// gt
disk[1632] <= 32'b010101_10011_00000_0000011001100101; 	// jf
disk[1633] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1634] <= 32'b111110_00000000000000010000101111; 	// jal
disk[1635] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1636] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1637] <= 32'b001111_11101_00101_0000000100011000; 	// lw
disk[1638] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1639] <= 32'b111100_00000000000000011001110100; 	// j
disk[1640] <= 32'b001111_11101_00101_0000000100100010; 	// lw
disk[1641] <= 32'b001111_11101_00110_0000000100100000; 	// lw
disk[1642] <= 32'b000000_00101_00110_10101_00000_001100; 	// eq
disk[1643] <= 32'b010101_10101_00000_0000011001110100; 	// jf
disk[1644] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1645] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[1646] <= 32'b000000_00111_10111_10110_00000_010000; 	// gt
disk[1647] <= 32'b010101_10110_00000_0000011001110100; 	// jf
disk[1648] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1649] <= 32'b111110_00000000000000001111111100; 	// jal
disk[1650] <= 32'b000010_11110_11110_0000000000000111; 	// subi
disk[1651] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1652] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1653] <= 32'b010010_11101_00101_0000000100100010; 	// sw
disk[1654] <= 32'b001111_11101_00110_0000000100100010; 	// lw
disk[1655] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1656] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[1657] <= 32'b111100_00000000000000010110000001; 	// j
disk[1658] <= 32'b111111_00000000000000000000000000; 	// halt

		// prog
disk[1700] <= 32'b111101_00000000000000000000010100;		// Jump to Main
disk[1701] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[1702] <= 32'b010010_11110_00001_1111111111111111; 	// sw
disk[1703] <= 32'b010000_00000_01111_0000000000000001; 	// li
disk[1704] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[1705] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[1706] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[1707] <= 32'b000000_00101_10001_10000_00000_010000; 	// gt
disk[1708] <= 32'b010101_10000_00000_0000000000010001; 	// jf
disk[1709] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[1710] <= 32'b000000_00110_00101_10010_00000_000010; 	// mul
disk[1711] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[1712] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[1713] <= 32'b000010_00101_10011_0000000000000001; 	// subi
disk[1714] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[1715] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[1716] <= 32'b111100_00000000000000000000000101; 	// j
disk[1717] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1718] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[1719] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[1720] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[1721] <= 32'b010000_00000_01111_0000000001011101; 	// li
disk[1722] <= 32'b010010_11110_01111_1111111111111110; 	// sw
disk[1723] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[1724] <= 32'b010010_11110_00101_1111111111111111; 	// sw
disk[1725] <= 32'b101000_00000000000000000000000000; 	// preIO
disk[1726] <= 32'b010011_00000_10000_0000000000000000; 	// in
disk[1727] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[1728] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1729] <= 32'b010000_00000_00010_0000000000000000; 	// li
disk[1730] <= 32'b010100_00000_00001_0000000000000000; 	// out
disk[1731] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[1732] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1733] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[1734] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[1735] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[1736] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1737] <= 32'b010010_11110_11111_1111111111111101; 	// sw
disk[1738] <= 32'b111110_00000000000000000000000001; 	// jal
disk[1739] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1740] <= 32'b001111_11110_11111_1111111111111101; 	// lw
disk[1741] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1742] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1743] <= 32'b010000_00000_00010_0000000000000010; 	// li
disk[1744] <= 32'b010100_00000_00001_0000000000000010; 	// out
disk[1745] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1746] <= 32'b011111_11001_00000_0000000000000000; 	// syscall


disk[1800] <= 32'b111101_00000000000000000000010010;		// Jump to Main
disk[1801] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[1802] <= 32'b010010_11110_00001_0000000000000000; 	// sw
disk[1803] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1804] <= 32'b000001_00101_01111_0000000000000001; 	// addi
disk[1805] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[1806] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1807] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1808] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[1809] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[1810] <= 32'b000001_00101_10000_0000000000000001; 	// addi
disk[1811] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[1812] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1813] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1814] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[1815] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[1816] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[1817] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[1818] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[1819] <= 32'b001110_11110_01111_0000000000000000; 	// mov
disk[1820] <= 32'b001110_01111_00001_0000000000000000; 	// mov
disk[1821] <= 32'b010000_00000_00010_0000000000000010; 	// li
disk[1822] <= 32'b010100_00000_00001_0000000000000010; 	// out
disk[1823] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[1824] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[1825] <= 32'b111110_00000000000000000000000001; 	// jal
disk[1826] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1827] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[1828] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1829] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[1830] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[1831] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1832] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[1833] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[1834] <= 32'b000001_00110_10000_0000000000000001; 	// addi
disk[1835] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[1836] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[1837] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1838] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[1839] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[1840] <= 32'b000001_00110_10001_0000000000000001; 	// addi
disk[1841] <= 32'b010010_11110_10001_0000000000000000; 	// sw
disk[1842] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[1843] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1844] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[1845] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[1846] <= 32'b000001_00110_10010_0000000000000001; 	// addi
disk[1847] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[1848] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[1849] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1850] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[1851] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[1852] <= 32'b000001_00110_10011_0000000000000001; 	// addi
disk[1853] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[1854] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[1855] <= 32'b010000_00000_00001_0000000000001011; 	// li
disk[1856] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[1857] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[1858] <= 32'b010000_00000_00001_0000000000001011; 	// li
disk[1859] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[1860] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[1861] <= 32'b001110_11110_10100_0000000000000000; 	// mov
disk[1862] <= 32'b001110_10100_00001_0000000000000000; 	// mov
disk[1863] <= 32'b010000_00000_00010_0000000000000010; 	// li
disk[1864] <= 32'b010100_00000_00001_0000000000000010; 	// out
disk[1865] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1866] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[1867] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[1868] <= 32'b000001_00110_10101_0000000000000001; 	// addi
disk[1869] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[1870] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[1871] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1872] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[1873] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[1874] <= 32'b000001_00110_10110_0000000000000001; 	// addi
disk[1875] <= 32'b010010_11110_10110_0000000000000000; 	// sw
disk[1876] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[1877] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1878] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[1879] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[1880] <= 32'b000001_00110_10111_0000000000000001; 	// addi
disk[1881] <= 32'b010010_11110_10111_0000000000000000; 	// sw
disk[1882] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[1883] <= 32'b010000_00000_00001_0000000000010110; 	// li
disk[1884] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[1885] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[1886] <= 32'b010000_00000_00001_0000000000010110; 	// li
disk[1887] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[1888] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[1889] <= 32'b001110_11110_01111_0000000000000000; 	// mov
disk[1890] <= 32'b001110_01111_00001_0000000000000000; 	// mov
disk[1891] <= 32'b010000_00000_00010_0000000000000010; 	// li
disk[1892] <= 32'b010100_00000_00001_0000000000000010; 	// out
disk[1893] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[1894] <= 32'b011111_11001_00000_0000000000000000; 	// syscall



	end
endmodule
