module disco_rigido (clk, we, addr, datain, dataout);
	input clk;										// clock
	input we;										// write enable
	input [31:0] addr;							// disk address
	input [31:0] datain;							// data in (to disk)
	
	output reg [31:0] dataout;					// data out (from disk)
	
	localparam DISK_SIZE = 2048;				// Tamanho do disco
	reg [31:0] disk [DISK_SIZE-1:0];			// disk cells
	
	always @ (posedge clk) begin
		if (we) disk[addr] <= datain;			// write disk
	end
	
	always @ (negedge clk) begin
		dataout <= disk[addr];
	end

	initial begin
		// SISTEMA OPERACIONAL

		
disk[0] <= 32'b111100_00000000000000001011111011;		// Jump to Main
disk[1] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[2] <= 32'b010010_11110_00001_0000000000000000; 	// sw
disk[3] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[4] <= 32'b001111_11101_00110_0000000001101101; 	// lw
disk[5] <= 32'b000000_00101_00110_01111_00000_000010; 	// mul
disk[6] <= 32'b001110_01111_00001_0000000000000000; 	// mov
disk[7] <= 32'b010010_00001_00000_0000000000000000; 	// sw
disk[8] <= 32'b010010_00001_00001_0000000000000001; 	// sw
disk[9] <= 32'b010010_00001_00010_0000000000000010; 	// sw
disk[10] <= 32'b010010_00001_00011_0000000000000011; 	// sw
disk[11] <= 32'b010010_00001_00100_0000000000000100; 	// sw
disk[12] <= 32'b010010_00001_00101_0000000000000101; 	// sw
disk[13] <= 32'b010010_00001_00110_0000000000000110; 	// sw
disk[14] <= 32'b010010_00001_00111_0000000000000111; 	// sw
disk[15] <= 32'b010010_00001_01000_0000000000001000; 	// sw
disk[16] <= 32'b010010_00001_01001_0000000000001001; 	// sw
disk[17] <= 32'b010010_00001_01010_0000000000001010; 	// sw
disk[18] <= 32'b010010_00001_01011_0000000000001011; 	// sw
disk[19] <= 32'b010010_00001_01100_0000000000001100; 	// sw
disk[20] <= 32'b010010_00001_01101_0000000000001101; 	// sw
disk[21] <= 32'b010010_00001_01110_0000000000001110; 	// sw
disk[22] <= 32'b010010_00001_01111_0000000000001111; 	// sw
disk[23] <= 32'b010010_00001_10000_0000000000010000; 	// sw
disk[24] <= 32'b010010_00001_10001_0000000000010001; 	// sw
disk[25] <= 32'b010010_00001_10010_0000000000010010; 	// sw
disk[26] <= 32'b010010_00001_10011_0000000000010011; 	// sw
disk[27] <= 32'b010010_00001_10100_0000000000010100; 	// sw
disk[28] <= 32'b010010_00001_10101_0000000000010101; 	// sw
disk[29] <= 32'b010010_00001_10110_0000000000010110; 	// sw
disk[30] <= 32'b010010_00001_10111_0000000000010111; 	// sw
disk[31] <= 32'b010010_00001_11000_0000000000011000; 	// sw
disk[32] <= 32'b010010_00001_11001_0000000000011001; 	// sw
disk[33] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[34] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[35] <= 32'b010010_11110_00001_0000000000000000; 	// sw
disk[36] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[37] <= 32'b001111_11101_00110_0000000001101101; 	// lw
disk[38] <= 32'b000000_00101_00110_01111_00000_000010; 	// mul
disk[39] <= 32'b001110_01111_00001_0000000000000000; 	// mov
disk[40] <= 32'b001111_00001_00000_0000000000000000; 	// lw
disk[41] <= 32'b001111_00001_00001_0000000000000001; 	// lw
disk[42] <= 32'b001111_00001_00010_0000000000000010; 	// lw
disk[43] <= 32'b001111_00001_00011_0000000000000011; 	// lw
disk[44] <= 32'b001111_00001_00100_0000000000000100; 	// lw
disk[45] <= 32'b001111_00001_00101_0000000000000101; 	// lw
disk[46] <= 32'b001111_00001_00110_0000000000000110; 	// lw
disk[47] <= 32'b001111_00001_00111_0000000000000111; 	// lw
disk[48] <= 32'b001111_00001_01000_0000000000001000; 	// lw
disk[49] <= 32'b001111_00001_01001_0000000000001001; 	// lw
disk[50] <= 32'b001111_00001_01010_0000000000001010; 	// lw
disk[51] <= 32'b001111_00001_01011_0000000000001011; 	// lw
disk[52] <= 32'b001111_00001_01100_0000000000001100; 	// lw
disk[53] <= 32'b001111_00001_01101_0000000000001101; 	// lw
disk[54] <= 32'b001111_00001_01110_0000000000001110; 	// lw
disk[55] <= 32'b001111_00001_01111_0000000000001111; 	// lw
disk[56] <= 32'b001111_00001_10000_0000000000010000; 	// lw
disk[57] <= 32'b001111_00001_10001_0000000000010001; 	// lw
disk[58] <= 32'b001111_00001_10010_0000000000010010; 	// lw
disk[59] <= 32'b001111_00001_10011_0000000000010011; 	// lw
disk[60] <= 32'b001111_00001_10100_0000000000010100; 	// lw
disk[61] <= 32'b001111_00001_10101_0000000000010101; 	// lw
disk[62] <= 32'b001111_00001_10110_0000000000010110; 	// lw
disk[63] <= 32'b001111_00001_10111_0000000000010111; 	// lw
disk[64] <= 32'b001111_00001_11000_0000000000011000; 	// lw
disk[65] <= 32'b001111_00001_11001_0000000000011001; 	// lw
disk[66] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[67] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[68] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[69] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[70] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[71] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[72] <= 32'b010110_00001_10000_0000000000000000; 	// ldk
disk[73] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[74] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[75] <= 32'b001101_00101_10001_0000000000011010; 	// srli
disk[76] <= 32'b001111_11101_00110_0000000010100010; 	// lw
disk[77] <= 32'b000000_10001_00110_10010_00000_001101; 	// ne
disk[78] <= 32'b010101_10010_00000_0000000001011000; 	// jf
disk[79] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[80] <= 32'b000001_00111_10011_0000000000000001; 	// addi
disk[81] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[82] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[83] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[84] <= 32'b010110_00001_10100_0000000000000000; 	// ldk
disk[85] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[86] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[87] <= 32'b111100_00000000000000000001001010; 	// j
disk[88] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[89] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[90] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[91] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[92] <= 32'b010010_11110_00001_1111111111111111; 	// sw
disk[93] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[94] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[95] <= 32'b000000_00101_10000_01111_00000_001100; 	// eq
disk[96] <= 32'b010101_01111_00000_0000000001100100; 	// jf
disk[97] <= 32'b010000_00000_10001_0000000000000001; 	// li
disk[98] <= 32'b001110_10001_11001_0000000000000000; 	// mov
disk[99] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[100] <= 32'b010000_00000_10010_0000000000000001; 	// li
disk[101] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[102] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[103] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[104] <= 32'b000000_00101_10100_10011_00000_010000; 	// gt
disk[105] <= 32'b010101_10011_00000_0000000001110010; 	// jf
disk[106] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[107] <= 32'b000011_00110_10101_0000000000000010; 	// muli
disk[108] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[109] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[110] <= 32'b000010_00101_10110_0000000000000001; 	// subi
disk[111] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[112] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[113] <= 32'b111100_00000000000000000001100110; 	// j
disk[114] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[115] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[116] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[117] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[118] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[119] <= 32'b010000_00000_00010_0000000000000000; 	// li
disk[120] <= 32'b010100_00000_00001_0000000000000000; 	// out
disk[121] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[122] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[123] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[124] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[125] <= 32'b010000_00000_00010_0000000000000010; 	// li
disk[126] <= 32'b010100_00000_00001_0000000000000010; 	// out
disk[127] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[128] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[129] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[130] <= 32'b010010_11101_01111_0000000001110011; 	// sw
disk[131] <= 32'b010000_00000_10000_0000000000000001; 	// li
disk[132] <= 32'b010010_11101_10000_0000000001110100; 	// sw
disk[133] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[134] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[135] <= 32'b010000_00000_01111_0000000000000001; 	// li
disk[136] <= 32'b010010_11101_01111_0000000000000000; 	// sw
disk[137] <= 32'b010000_00000_10000_0000000000000010; 	// li
disk[138] <= 32'b010010_11101_10000_0000000000000001; 	// sw
disk[139] <= 32'b010000_00000_10001_0000000000000011; 	// li
disk[140] <= 32'b010010_11101_10001_0000000000000010; 	// sw
disk[141] <= 32'b010000_00000_10010_0000000110010100; 	// li
disk[142] <= 32'b010010_11101_10010_0000000000000011; 	// sw
disk[143] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[144] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[145] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[146] <= 32'b010000_00000_10101_0000000000001010; 	// li
disk[147] <= 32'b000000_00101_10101_10100_00000_001110; 	// lt
disk[148] <= 32'b010101_10100_00000_0000000010101001; 	// jf
disk[149] <= 32'b010001_11101_00110_0000000000000100; 	// la
disk[150] <= 32'b000000_00110_00101_10110_00000_000000; 	// add
disk[151] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[152] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[153] <= 32'b010001_11101_00111_0000000000001110; 	// la
disk[154] <= 32'b000000_00111_00101_11000_00000_000000; 	// add
disk[155] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[156] <= 32'b010010_11000_01111_0000000000000000; 	// sw
disk[157] <= 32'b010001_11101_01000_0000000000011000; 	// la
disk[158] <= 32'b000000_01000_00101_10000_00000_000000; 	// add
disk[159] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[160] <= 32'b010010_10000_10001_0000000000000000; 	// sw
disk[161] <= 32'b010001_11101_01001_0000000000100010; 	// la
disk[162] <= 32'b000000_01001_00101_10010_00000_000000; 	// add
disk[163] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[164] <= 32'b010010_10010_10011_0000000000000000; 	// sw
disk[165] <= 32'b000001_00101_10100_0000000000000001; 	// addi
disk[166] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[167] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[168] <= 32'b111100_00000000000000000010010001; 	// j
disk[169] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[170] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[171] <= 32'b010000_00000_01111_0000000000100000; 	// li
disk[172] <= 32'b010010_11101_01111_0000000001101101; 	// sw
disk[173] <= 32'b010000_00000_10000_0000000001000000; 	// li
disk[174] <= 32'b010010_11101_10000_0000000001101110; 	// sw
disk[175] <= 32'b010000_00000_10001_0000000001100100; 	// li
disk[176] <= 32'b010010_11101_10001_0000000001101111; 	// sw
disk[177] <= 32'b010000_00000_10010_0000000000001010; 	// li
disk[178] <= 32'b010010_11101_10010_0000000001110000; 	// sw
disk[179] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[180] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[181] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[182] <= 32'b010010_11101_01111_0000000010100011; 	// sw
disk[183] <= 32'b010000_00000_10000_0000000000000001; 	// li
disk[184] <= 32'b010010_11101_10000_0000000010100100; 	// sw
disk[185] <= 32'b010000_00000_10001_0000000000000010; 	// li
disk[186] <= 32'b010010_11101_10001_0000000010100101; 	// sw
disk[187] <= 32'b010000_00000_10010_0000000000000011; 	// li
disk[188] <= 32'b010010_11101_10010_0000000010100110; 	// sw
disk[189] <= 32'b010000_00000_10011_0000000000000100; 	// li
disk[190] <= 32'b010010_11101_10011_0000000010100111; 	// sw
disk[191] <= 32'b010000_00000_10100_0000000000000101; 	// li
disk[192] <= 32'b010010_11101_10100_0000000010101000; 	// sw
disk[193] <= 32'b010000_00000_10101_0000000000001010; 	// li
disk[194] <= 32'b010010_11101_10101_0000000010101001; 	// sw
disk[195] <= 32'b001111_11101_00101_0000000010100011; 	// lw
disk[196] <= 32'b010010_11101_00101_0000000010101010; 	// sw
disk[197] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[198] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[199] <= 32'b010000_00000_01111_0000011111111111; 	// li
disk[200] <= 32'b010010_11101_01111_0000000001110010; 	// sw
disk[201] <= 32'b010000_00000_10000_0000000000011111; 	// li
disk[202] <= 32'b010010_11101_10000_0000000010100000; 	// sw
disk[203] <= 32'b010000_00000_10001_0000000000111101; 	// li
disk[204] <= 32'b010010_11101_10001_0000000010100001; 	// sw
disk[205] <= 32'b010000_00000_10010_0000000000111111; 	// li
disk[206] <= 32'b010010_11101_10010_0000000010100010; 	// sw
disk[207] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[208] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[209] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[210] <= 32'b010010_11110_01111_1111111111111110; 	// sw
disk[211] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[212] <= 32'b001111_11101_00110_0000000001101110; 	// lw
disk[213] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[214] <= 32'b010101_10000_00000_0000000011011111; 	// jf
disk[215] <= 32'b010001_11101_00111_0000000000101101; 	// la
disk[216] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[217] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[218] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[219] <= 32'b000001_00101_10011_0000000000000001; 	// addi
disk[220] <= 32'b010010_11110_10011_1111111111111110; 	// sw
disk[221] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[222] <= 32'b111100_00000000000000000011010011; 	// j
disk[223] <= 32'b010010_11110_11111_1111111111111101; 	// sw
disk[224] <= 32'b111110_00000000000000000001000011; 	// jal
disk[225] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[226] <= 32'b001111_11110_11111_1111111111111101; 	// lw
disk[227] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[228] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[229] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[230] <= 32'b000001_00110_10100_0000000000000001; 	// addi
disk[231] <= 32'b010010_11101_10100_0000000001110001; 	// sw
disk[232] <= 32'b001111_11101_00111_0000000001101101; 	// lw
disk[233] <= 32'b000000_00110_00111_10101_00000_000011; 	// div
disk[234] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[235] <= 32'b000000_00110_00111_10110_00000_000100; 	// mod
disk[236] <= 32'b010000_00000_11000_0000000000000000; 	// li
disk[237] <= 32'b000000_10110_11000_10111_00000_010000; 	// gt
disk[238] <= 32'b010101_10111_00000_0000000011110011; 	// jf
disk[239] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[240] <= 32'b000001_01000_01111_0000000000000001; 	// addi
disk[241] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[242] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[243] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[244] <= 32'b010010_11110_10000_1111111111111110; 	// sw
disk[245] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[246] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[247] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[248] <= 32'b010101_10001_00000_0000000100000001; 	// jf
disk[249] <= 32'b010001_11101_00111_0000000000101101; 	// la
disk[250] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
disk[251] <= 32'b010000_00000_10011_0000000000000001; 	// li
disk[252] <= 32'b010010_10010_10011_0000000000000000; 	// sw
disk[253] <= 32'b000001_00101_10100_0000000000000001; 	// addi
disk[254] <= 32'b010010_11110_10100_1111111111111110; 	// sw
disk[255] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[256] <= 32'b111100_00000000000000000011110101; 	// j
disk[257] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[258] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[259] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[260] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[261] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[262] <= 32'b001111_11101_00110_0000000001110000; 	// lw
disk[263] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[264] <= 32'b010101_10000_00000_0000000100011101; 	// jf
disk[265] <= 32'b010001_11101_00111_0000000001111000; 	// la
disk[266] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[267] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[268] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[269] <= 32'b010001_11101_01000_0000000010000010; 	// la
disk[270] <= 32'b000000_01000_00101_10011_00000_000000; 	// add
disk[271] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[272] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[273] <= 32'b010001_11101_01001_0000000010001100; 	// la
disk[274] <= 32'b000000_01001_00101_10101_00000_000000; 	// add
disk[275] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[276] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[277] <= 32'b010001_11101_01010_0000000010010110; 	// la
disk[278] <= 32'b000000_01010_00101_10111_00000_000000; 	// add
disk[279] <= 32'b010000_00000_11000_0000000000000000; 	// li
disk[280] <= 32'b010010_10111_11000_0000000000000000; 	// sw
disk[281] <= 32'b000001_00101_01111_0000000000000001; 	// addi
disk[282] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[283] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[284] <= 32'b111100_00000000000000000100000101; 	// j
disk[285] <= 32'b001111_11101_00101_0000000001110001; 	// lw
disk[286] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[287] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[288] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[289] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[290] <= 32'b001111_11101_00110_0000000001110010; 	// lw
disk[291] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[292] <= 32'b010101_10001_00000_0000000100111101; 	// jf
disk[293] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[294] <= 32'b010110_00001_10010_0000000000000000; 	// ldk
disk[295] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[296] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[297] <= 32'b001101_00111_10011_0000000000011010; 	// srli
disk[298] <= 32'b001111_11101_01000_0000000010100001; 	// lw
disk[299] <= 32'b000000_10011_01000_10100_00000_001100; 	// eq
disk[300] <= 32'b010101_10100_00000_0000000100111000; 	// jf
disk[301] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[302] <= 32'b000001_01001_10101_0000000000000001; 	// addi
disk[303] <= 32'b010001_11101_01010_0000000001111000; 	// la
disk[304] <= 32'b000000_01010_01001_10110_00000_000000; 	// add
disk[305] <= 32'b010010_10110_10101_0000000000000000; 	// sw
disk[306] <= 32'b010001_11101_01011_0000000010000010; 	// la
disk[307] <= 32'b000000_01011_01001_10111_00000_000000; 	// add
disk[308] <= 32'b010010_10111_00101_0000000000000000; 	// sw
disk[309] <= 32'b000001_01001_11000_0000000000000001; 	// addi
disk[310] <= 32'b010010_11110_11000_1111111111111111; 	// sw
disk[311] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[312] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[313] <= 32'b000001_00101_01111_0000000000000001; 	// addi
disk[314] <= 32'b010010_11110_01111_1111111111111110; 	// sw
disk[315] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[316] <= 32'b111100_00000000000000000100100001; 	// j
disk[317] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[318] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[319] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[320] <= 32'b111110_00000000000000000010000110; 	// jal
disk[321] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[322] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[323] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[324] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[325] <= 32'b111110_00000000000000000010101010; 	// jal
disk[326] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[327] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[328] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[329] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[330] <= 32'b111110_00000000000000000010110100; 	// jal
disk[331] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[332] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[333] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[334] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[335] <= 32'b111110_00000000000000000011000110; 	// jal
disk[336] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[337] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[338] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[339] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[340] <= 32'b111110_00000000000000000011010000; 	// jal
disk[341] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[342] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[343] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[344] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[345] <= 32'b111110_00000000000000000100000010; 	// jal
disk[346] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[347] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[348] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[349] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[350] <= 32'b000001_11110_11110_0000000000000110; 	// addi
disk[351] <= 32'b010010_11110_00001_1111111111111101; 	// sw
disk[352] <= 32'b001111_11110_00101_1111111111111101; 	// lw
disk[353] <= 32'b001111_11101_00110_0000000001101101; 	// lw
disk[354] <= 32'b000000_00101_00110_01111_00000_000011; 	// div
disk[355] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[356] <= 32'b000000_00101_00110_10000_00000_000100; 	// mod
disk[357] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[358] <= 32'b000000_10000_10010_10001_00000_010000; 	// gt
disk[359] <= 32'b010101_10001_00000_0000000101101100; 	// jf
disk[360] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[361] <= 32'b000001_00111_10011_0000000000000001; 	// addi
disk[362] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[363] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[364] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[365] <= 32'b010010_11110_10100_1111111111111110; 	// sw
disk[366] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[367] <= 32'b001111_11101_00110_0000000001101110; 	// lw
disk[368] <= 32'b000000_00101_00110_10101_00000_001110; 	// lt
disk[369] <= 32'b010101_10101_00000_0000000110010001; 	// jf
disk[370] <= 32'b010001_11101_00111_0000000000101101; 	// la
disk[371] <= 32'b000000_00111_00101_10110_00000_000000; 	// add
disk[372] <= 32'b001111_10110_10110_0000000000000000; 	// lw
disk[373] <= 32'b010000_00000_11000_0000000000000000; 	// li
disk[374] <= 32'b000000_10110_11000_10111_00000_001100; 	// eq
disk[375] <= 32'b010101_10111_00000_0000000110001100; 	// jf
disk[376] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[377] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[378] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[379] <= 32'b000000_00101_10000_01111_00000_001101; 	// ne
disk[380] <= 32'b010101_01111_00000_0000000110001001; 	// jf
disk[381] <= 32'b010001_11101_00110_0000000000101101; 	// la
disk[382] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[383] <= 32'b000000_00110_00111_10001_00000_000000; 	// add
disk[384] <= 32'b010000_00000_10010_0000000000000001; 	// li
disk[385] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[386] <= 32'b000010_00101_10011_0000000000000001; 	// subi
disk[387] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[388] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[389] <= 32'b000001_00111_10100_0000000000000001; 	// addi
disk[390] <= 32'b010010_11110_10100_1111111111111110; 	// sw
disk[391] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[392] <= 32'b111100_00000000000000000101111001; 	// j
disk[393] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[394] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[395] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[396] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[397] <= 32'b000001_00101_10101_0000000000000001; 	// addi
disk[398] <= 32'b010010_11110_10101_1111111111111110; 	// sw
disk[399] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[400] <= 32'b111100_00000000000000000101101110; 	// j
disk[401] <= 32'b001111_11101_00101_0000000001101111; 	// lw
disk[402] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[403] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[404] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[405] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[406] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[407] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[408] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[409] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[410] <= 32'b001111_11101_00110_0000000001110000; 	// lw
disk[411] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[412] <= 32'b010101_10001_00000_0000000110110010; 	// jf
disk[413] <= 32'b010001_11101_00111_0000000010001100; 	// la
disk[414] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
disk[415] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[416] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[417] <= 32'b000000_10010_10100_10011_00000_001101; 	// ne
disk[418] <= 32'b010101_10011_00000_0000000110101101; 	// jf
disk[419] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[420] <= 32'b010010_11110_11111_1111111111111110; 	// sw
disk[421] <= 32'b111110_00000000000000000001011011; 	// jal
disk[422] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[423] <= 32'b001111_11110_11111_1111111111111110; 	// lw
disk[424] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[425] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[426] <= 32'b000000_00110_00101_10101_00000_000000; 	// add
disk[427] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[428] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[429] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[430] <= 32'b000001_00101_10110_0000000000000001; 	// addi
disk[431] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[432] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[433] <= 32'b111100_00000000000000000110011001; 	// j
disk[434] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[435] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[436] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[437] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[438] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[439] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[440] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[441] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[442] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[443] <= 32'b001111_11101_00110_0000000001110000; 	// lw
disk[444] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[445] <= 32'b010101_10001_00000_0000000111010011; 	// jf
disk[446] <= 32'b010001_11101_00111_0000000001111000; 	// la
disk[447] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
disk[448] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[449] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[450] <= 32'b000000_10010_10100_10011_00000_001101; 	// ne
disk[451] <= 32'b010101_10011_00000_0000000111001110; 	// jf
disk[452] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[453] <= 32'b010010_11110_11111_1111111111111110; 	// sw
disk[454] <= 32'b111110_00000000000000000001011011; 	// jal
disk[455] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[456] <= 32'b001111_11110_11111_1111111111111110; 	// lw
disk[457] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[458] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[459] <= 32'b000000_00110_00101_10101_00000_000000; 	// add
disk[460] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[461] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[462] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[463] <= 32'b000001_00101_10110_0000000000000001; 	// addi
disk[464] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[465] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[466] <= 32'b111100_00000000000000000110111010; 	// j
disk[467] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[468] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[469] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[470] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[471] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[472] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[473] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[474] <= 32'b001111_11101_00110_0000000001110000; 	// lw
disk[475] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[476] <= 32'b010101_10000_00000_0000000111101010; 	// jf
disk[477] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[478] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[479] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[480] <= 32'b001111_11101_01000_0000000000000010; 	// lw
disk[481] <= 32'b000000_10001_01000_10010_00000_001100; 	// eq
disk[482] <= 32'b010101_10010_00000_0000000111100101; 	// jf
disk[483] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[484] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[485] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[486] <= 32'b000001_00101_10011_0000000000000001; 	// addi
disk[487] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[488] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[489] <= 32'b111100_00000000000000000111011001; 	// j
disk[490] <= 32'b001111_11101_00101_0000000000000011; 	// lw
disk[491] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[492] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[493] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[494] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[495] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[496] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[497] <= 32'b001111_11101_00110_0000000001110000; 	// lw
disk[498] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[499] <= 32'b010101_10000_00000_0000001000000001; 	// jf
disk[500] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[501] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[502] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[503] <= 32'b001111_11101_01000_0000000000000001; 	// lw
disk[504] <= 32'b000000_10001_01000_10010_00000_001100; 	// eq
disk[505] <= 32'b010101_10010_00000_0000000111111100; 	// jf
disk[506] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[507] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[508] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[509] <= 32'b000001_00101_10011_0000000000000001; 	// addi
disk[510] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[511] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[512] <= 32'b111100_00000000000000000111110000; 	// j
disk[513] <= 32'b001111_11101_00101_0000000000000011; 	// lw
disk[514] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[515] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[516] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[517] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[518] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[519] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[520] <= 32'b001111_11101_00110_0000000001110000; 	// lw
disk[521] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[522] <= 32'b010101_10000_00000_0000001000011010; 	// jf
disk[523] <= 32'b010001_11101_00111_0000000010001100; 	// la
disk[524] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[525] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[526] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[527] <= 32'b000000_10001_10011_10010_00000_001101; 	// ne
disk[528] <= 32'b010101_10010_00000_0000001000010101; 	// jf
disk[529] <= 32'b010001_11101_01000_0000000000000100; 	// la
disk[530] <= 32'b000000_01000_00101_10100_00000_000000; 	// add
disk[531] <= 32'b001111_11101_01001_0000000000000001; 	// lw
disk[532] <= 32'b010010_10100_01001_0000000000000000; 	// sw
disk[533] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[534] <= 32'b000001_00101_10101_0000000000000001; 	// addi
disk[535] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[536] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[537] <= 32'b111100_00000000000000001000000111; 	// j
disk[538] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[539] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[540] <= 32'b010010_11110_00001_1111111111111110; 	// sw
disk[541] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[542] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[543] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[544] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[545] <= 32'b010110_00001_01111_0000000000000000; 	// ldk
disk[546] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[547] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[548] <= 32'b001101_00101_10000_0000000000011010; 	// srli
disk[549] <= 32'b001111_11101_00110_0000000010100000; 	// lw
disk[550] <= 32'b000000_10000_00110_10001_00000_001101; 	// ne
disk[551] <= 32'b010101_10001_00000_0000001000110001; 	// jf
disk[552] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[553] <= 32'b000001_00111_10010_0000000000000001; 	// addi
disk[554] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[555] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[556] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[557] <= 32'b010110_00001_10011_0000000000000000; 	// ldk
disk[558] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[559] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[560] <= 32'b111100_00000000000000001000100011; 	// j
disk[561] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[562] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[563] <= 32'b000000_00101_00110_10100_00000_000001; 	// sub
disk[564] <= 32'b001110_10100_11001_0000000000000000; 	// mov
disk[565] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[566] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[567] <= 32'b010010_11110_00001_0000000000000001; 	// sw
disk[568] <= 32'b001111_11110_00101_0000000000000001; 	// lw
disk[569] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[570] <= 32'b010010_11110_01111_0000000000000001; 	// sw
disk[571] <= 32'b001111_11110_00101_0000000000000001; 	// lw
disk[572] <= 32'b010001_11101_00110_0000000010000010; 	// la
disk[573] <= 32'b000000_00110_00101_10000_00000_000000; 	// add
disk[574] <= 32'b001111_10000_10000_0000000000000000; 	// lw
disk[575] <= 32'b010010_11110_10000_0000000000000111; 	// sw
disk[576] <= 32'b010001_11101_00111_0000000001111000; 	// la
disk[577] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[578] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[579] <= 32'b010010_11110_10001_0000000000001000; 	// sw
disk[580] <= 32'b001111_11110_01000_0000000000000111; 	// lw
disk[581] <= 32'b010010_11110_01000_0000000000000010; 	// sw
disk[582] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[583] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[584] <= 32'b111110_00000000000000001000011011; 	// jal
disk[585] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[586] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[587] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[588] <= 32'b010010_11110_00101_0000000000000110; 	// sw
disk[589] <= 32'b001111_11110_00110_0000000000000110; 	// lw
disk[590] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[591] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[592] <= 32'b111110_00000000000000000101011110; 	// jal
disk[593] <= 32'b000010_11110_11110_0000000000000110; 	// subi
disk[594] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[595] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[596] <= 32'b010010_11110_00101_0000000000000101; 	// sw
disk[597] <= 32'b001111_11101_00110_0000000001101101; 	// lw
disk[598] <= 32'b001111_11110_00111_0000000000000101; 	// lw
disk[599] <= 32'b000000_00110_00111_10010_00000_000010; 	// mul
disk[600] <= 32'b010010_11110_10010_0000000000000011; 	// sw
disk[601] <= 32'b001111_11110_01000_0000000000000010; 	// lw
disk[602] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[603] <= 32'b010110_00001_10011_0000000000000000; 	// ldk
disk[604] <= 32'b010010_11110_10011_0000000000000100; 	// sw
disk[605] <= 32'b001111_11110_00101_0000000000000100; 	// lw
disk[606] <= 32'b001101_00101_10100_0000000000011010; 	// srli
disk[607] <= 32'b001111_11101_00110_0000000010100000; 	// lw
disk[608] <= 32'b000000_10100_00110_10101_00000_001101; 	// ne
disk[609] <= 32'b010101_10101_00000_0000001001110010; 	// jf
disk[610] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[611] <= 32'b001111_11110_00111_0000000000000011; 	// lw
disk[612] <= 32'b001110_00111_00010_0000000000000000; 	// mov
disk[613] <= 32'b011001_00010_00001_0000000000000000; 	// sim
disk[614] <= 32'b001111_11110_01000_0000000000000010; 	// lw
disk[615] <= 32'b000001_01000_10110_0000000000000001; 	// addi
disk[616] <= 32'b010010_11110_10110_0000000000000010; 	// sw
disk[617] <= 32'b001111_11110_01000_0000000000000010; 	// lw
disk[618] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[619] <= 32'b010110_00001_10111_0000000000000000; 	// ldk
disk[620] <= 32'b010010_11110_10111_0000000000000100; 	// sw
disk[621] <= 32'b001111_11110_00101_0000000000000100; 	// lw
disk[622] <= 32'b000001_00111_11000_0000000000000001; 	// addi
disk[623] <= 32'b010010_11110_11000_0000000000000011; 	// sw
disk[624] <= 32'b001111_11110_00111_0000000000000011; 	// lw
disk[625] <= 32'b111100_00000000000000001001011101; 	// j
disk[626] <= 32'b001111_11110_00101_0000000000000100; 	// lw
disk[627] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[628] <= 32'b001111_11110_00110_0000000000000011; 	// lw
disk[629] <= 32'b001110_00110_00010_0000000000000000; 	// mov
disk[630] <= 32'b011001_00010_00001_0000000000000000; 	// sim
disk[631] <= 32'b001111_11110_00111_0000000000001000; 	// lw
disk[632] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[633] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
disk[634] <= 32'b001111_11101_01000_0000000001101101; 	// lw
disk[635] <= 32'b001111_11110_01001_0000000000000101; 	// lw
disk[636] <= 32'b000000_01000_01001_01111_00000_000010; 	// mul
disk[637] <= 32'b001110_01111_00001_0000000000000000; 	// mov
disk[638] <= 32'b011010_00000_00001_0000000000000000; 	// mmuLowerIM
disk[639] <= 32'b010001_11101_01010_0000000010001100; 	// la
disk[640] <= 32'b001111_11110_01011_0000000000000001; 	// lw
disk[641] <= 32'b000000_01010_01011_10000_00000_000000; 	// add
disk[642] <= 32'b010010_10000_00111_0000000000000000; 	// sw
disk[643] <= 32'b010001_11101_01100_0000000010010110; 	// la
disk[644] <= 32'b000000_01100_01011_10001_00000_000000; 	// add
disk[645] <= 32'b001111_11110_01101_0000000000000111; 	// lw
disk[646] <= 32'b010010_10001_01101_0000000000000000; 	// sw
disk[647] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[648] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[649] <= 32'b010010_11110_00001_0000000000000000; 	// sw
disk[650] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[651] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[652] <= 32'b100100_00000_00001_0000000000000000; 	// lcdCurr
disk[653] <= 32'b001111_11101_00110_0000000010101001; 	// lw
disk[654] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[655] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[656] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[657] <= 32'b001111_11101_01000_0000000000101100; 	// lw
disk[658] <= 32'b000000_00111_01000_01111_00000_000000; 	// add
disk[659] <= 32'b001111_11101_01001_0000000000000000; 	// lw
disk[660] <= 32'b010010_01111_01001_0000000000000000; 	// sw
disk[661] <= 32'b010001_11101_01010_0000000000001110; 	// la
disk[662] <= 32'b000000_01010_01000_10000_00000_000000; 	// add
disk[663] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[664] <= 32'b010010_10000_10001_0000000000000000; 	// sw
disk[665] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[666] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
disk[667] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[668] <= 32'b100000_00000000000000000000000000; 	// exec
disk[669] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[670] <= 32'b010001_11101_00101_0000000000000100; 	// la
disk[671] <= 32'b001111_11101_00110_0000000000101100; 	// lw
disk[672] <= 32'b000000_00101_00110_10010_00000_000000; 	// add
disk[673] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[674] <= 32'b010010_10010_10011_0000000000000000; 	// sw
disk[675] <= 32'b010001_11101_00111_0000000000001110; 	// la
disk[676] <= 32'b000000_00111_00110_10100_00000_000000; 	// add
disk[677] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[678] <= 32'b010010_10100_10101_0000000000000000; 	// sw
disk[679] <= 32'b001111_11101_01000_0000000010100011; 	// lw
disk[680] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[681] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[682] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[683] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[684] <= 32'b010010_11110_00001_0000000000000000; 	// sw
disk[685] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[686] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[687] <= 32'b100100_00000_00001_0000000000000000; 	// lcdCurr
disk[688] <= 32'b001111_11101_00110_0000000010101001; 	// lw
disk[689] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[690] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[691] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[692] <= 32'b001111_11101_01000_0000000000101100; 	// lw
disk[693] <= 32'b000000_00111_01000_01111_00000_000000; 	// add
disk[694] <= 32'b001111_11101_01001_0000000000000000; 	// lw
disk[695] <= 32'b010010_01111_01001_0000000000000000; 	// sw
disk[696] <= 32'b000001_01000_10000_0000000000000001; 	// addi
disk[697] <= 32'b001110_10000_00001_0000000000000000; 	// mov
disk[698] <= 32'b010001_11101_01010_0000000000001110; 	// la
disk[699] <= 32'b000000_01010_01000_10001_00000_000000; 	// add
disk[700] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[701] <= 32'b001110_10001_00010_0000000000000000; 	// mov
disk[702] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
disk[703] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[704] <= 32'b001110_11100_11110_0000000000000000; 	// mov
disk[705] <= 32'b001110_11011_11101_0000000000000000; 	// mov
disk[706] <= 32'b100001_00010_00000_0000000000000000; 	// execAgain
disk[707] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[708] <= 32'b010001_11101_00101_0000000000000100; 	// la
disk[709] <= 32'b001111_11101_00110_0000000000101100; 	// lw
disk[710] <= 32'b000000_00101_00110_10010_00000_000000; 	// add
disk[711] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[712] <= 32'b010010_10010_10011_0000000000000000; 	// sw
disk[713] <= 32'b010001_11101_00111_0000000000001110; 	// la
disk[714] <= 32'b000000_00111_00110_10100_00000_000000; 	// add
disk[715] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[716] <= 32'b010010_10100_10101_0000000000000000; 	// sw
disk[717] <= 32'b001111_11101_01000_0000000010100011; 	// lw
disk[718] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[719] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[720] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[721] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[722] <= 32'b010010_11110_00001_0000000000000000; 	// sw
disk[723] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[724] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[725] <= 32'b010010_11101_01111_0000000000101100; 	// sw
disk[726] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[727] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[728] <= 32'b111110_00000000000000001010001000; 	// jal
disk[729] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[730] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[731] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[732] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[733] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[734] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[735] <= 32'b111110_00000000000000001000000100; 	// jal
disk[736] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[737] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[738] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[739] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[740] <= 32'b111110_00000000000000000111101101; 	// jal
disk[741] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[742] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[743] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[744] <= 32'b001111_11101_00110_0000000000000011; 	// lw
disk[745] <= 32'b000000_00101_00110_01111_00000_001101; 	// ne
disk[746] <= 32'b010101_01111_00000_0000001011111010; 	// jf
disk[747] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[748] <= 32'b111110_00000000000000000111101101; 	// jal
disk[749] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[750] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[751] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[752] <= 32'b010010_11101_00101_0000000000101100; 	// sw
disk[753] <= 32'b001111_11101_00110_0000000000101100; 	// lw
disk[754] <= 32'b000001_00110_10000_0000000000000001; 	// addi
disk[755] <= 32'b001110_10000_00001_0000000000000000; 	// mov
disk[756] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[757] <= 32'b111110_00000000000000001010001000; 	// jal
disk[758] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[759] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[760] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[761] <= 32'b111100_00000000000000001011100011; 	// j
disk[762] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[763] <= 32'b001110_11110_11100_0000000000000000; 	// mov
disk[764] <= 32'b001110_11101_11011_0000000000000000; 	// mov
disk[765] <= 32'b010000_00000_00000_0000000000000000; 	// li
disk[766] <= 32'b010000_00000_11110_0000000000000000; 	// li
disk[767] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[768] <= 32'b000001_11110_11110_0000000010101111; 	// addi
disk[769] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[770] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[771] <= 32'b000000_00101_10000_01111_00000_001100; 	// eq
disk[772] <= 32'b010101_01111_00000_0000001100001110; 	// jf
disk[773] <= 32'b111110_00000000000000000100111110; 	// jal
disk[774] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[775] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[776] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[777] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[778] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[779] <= 32'b010000_00000_10001_0000000000000001; 	// li
disk[780] <= 32'b010010_11110_10001_0000000000000000; 	// sw
disk[781] <= 32'b100110_00000_00000_0000000000000000; 	// cic
disk[782] <= 32'b100101_00000_10010_0000000000000000; 	// gic
disk[783] <= 32'b010010_11110_10010_1111111111111111; 	// sw
disk[784] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[785] <= 32'b010000_00000_10100_0000000000000001; 	// li
disk[786] <= 32'b000000_00101_10100_10011_00000_001100; 	// eq
disk[787] <= 32'b010101_10011_00000_0000001100101001; 	// jf
disk[788] <= 32'b010001_11101_00110_0000000000000100; 	// la
disk[789] <= 32'b001111_11101_00111_0000000000101100; 	// lw
disk[790] <= 32'b000000_00110_00111_10101_00000_000000; 	// add
disk[791] <= 32'b001111_11101_01000_0000000000000010; 	// lw
disk[792] <= 32'b010010_10101_01000_0000000000000000; 	// sw
disk[793] <= 32'b100111_00000_10110_0000000000000000; 	// gip
disk[794] <= 32'b000001_10110_10111_0000000000000001; 	// addi
disk[795] <= 32'b010001_11101_01001_0000000000001110; 	// la
disk[796] <= 32'b000000_01001_00111_11000_00000_000000; 	// add
disk[797] <= 32'b010010_11000_10111_0000000000000000; 	// sw
disk[798] <= 32'b100110_00000_00000_0000000000000000; 	// cic
disk[799] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[800] <= 32'b111110_00000000000000001010101011; 	// jal
disk[801] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[802] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[803] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[804] <= 32'b010000_00000_11110_0000000010101111; 	// li
disk[805] <= 32'b001110_11100_01111_0000000000000000; 	// mov
disk[806] <= 32'b001110_01111_00001_0000000000000000; 	// mov
disk[807] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[808] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[809] <= 32'b010000_00000_10000_0000000000000001; 	// li
disk[810] <= 32'b010101_10000_00000_0000001111000010; 	// jf
disk[811] <= 32'b010011_00000_10001_0000000000000000; 	// in
disk[812] <= 32'b010010_11110_10001_1111111111111110; 	// sw
disk[813] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[814] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[815] <= 32'b010000_00000_00010_0000000000000000; 	// li
disk[816] <= 32'b010100_00000_00001_0000000000000000; 	// out
disk[817] <= 32'b001111_11101_00110_0000000010101010; 	// lw
disk[818] <= 32'b001111_11101_00111_0000000010100011; 	// lw
disk[819] <= 32'b000000_00110_00111_10010_00000_001100; 	// eq
disk[820] <= 32'b010101_10010_00000_0000001101001101; 	// jf
disk[821] <= 32'b010000_00000_10100_0000000000000100; 	// li
disk[822] <= 32'b000000_00101_10100_10011_00000_010000; 	// gt
disk[823] <= 32'b010101_10011_00000_0000001100111011; 	// jf
disk[824] <= 32'b010010_11110_00111_1111111111111110; 	// sw
disk[825] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[826] <= 32'b111100_00000000000000001101001100; 	// j
disk[827] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[828] <= 32'b010000_00000_10110_0000000000000100; 	// li
disk[829] <= 32'b000000_00101_10110_10101_00000_001100; 	// eq
disk[830] <= 32'b010101_10101_00000_0000001101000101; 	// jf
disk[831] <= 32'b111110_00000000000000000001110101; 	// jal
disk[832] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[833] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[834] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[835] <= 32'b010010_11110_00110_1111111111111110; 	// sw
disk[836] <= 32'b111100_00000000000000001101001100; 	// j
disk[837] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[838] <= 32'b010000_00000_11000_0000000000000001; 	// li
disk[839] <= 32'b000000_00101_11000_10111_00000_001110; 	// lt
disk[840] <= 32'b010101_10111_00000_0000001101001100; 	// jf
disk[841] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[842] <= 32'b010010_11110_00110_1111111111111110; 	// sw
disk[843] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[844] <= 32'b111100_00000000000000001110111100; 	// j
disk[845] <= 32'b001111_11101_00101_0000000010101010; 	// lw
disk[846] <= 32'b001111_11101_00110_0000000010100100; 	// lw
disk[847] <= 32'b000000_00101_00110_01111_00000_001100; 	// eq
disk[848] <= 32'b010101_01111_00000_0000001101100001; 	// jf
disk[849] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[850] <= 32'b010000_00000_10001_0000000000000011; 	// li
disk[851] <= 32'b000000_00111_10001_10000_00000_010000; 	// gt
disk[852] <= 32'b010101_10000_00000_0000001101011001; 	// jf
disk[853] <= 32'b001111_11101_01000_0000000010100011; 	// lw
disk[854] <= 32'b010010_11110_01000_1111111111111110; 	// sw
disk[855] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[856] <= 32'b111100_00000000000000001101100000; 	// j
disk[857] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[858] <= 32'b010000_00000_10011_0000000000000001; 	// li
disk[859] <= 32'b000000_00101_10011_10010_00000_001110; 	// lt
disk[860] <= 32'b010101_10010_00000_0000001101100000; 	// jf
disk[861] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[862] <= 32'b010010_11110_00110_1111111111111110; 	// sw
disk[863] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[864] <= 32'b111100_00000000000000001110111100; 	// j
disk[865] <= 32'b001111_11101_00101_0000000010101010; 	// lw
disk[866] <= 32'b001111_11101_00110_0000000010100101; 	// lw
disk[867] <= 32'b000000_00101_00110_10100_00000_001100; 	// eq
disk[868] <= 32'b010101_10100_00000_0000001110000010; 	// jf
disk[869] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[870] <= 32'b010000_00000_10110_0000000000000001; 	// li
disk[871] <= 32'b000000_00111_10110_10101_00000_001100; 	// eq
disk[872] <= 32'b010101_10101_00000_0000001101110010; 	// jf
disk[873] <= 32'b001111_11101_01000_0000000010100111; 	// lw
disk[874] <= 32'b010010_11110_01000_1111111111111110; 	// sw
disk[875] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[876] <= 32'b111110_00000000000000000110110101; 	// jal
disk[877] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[878] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[879] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[880] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[881] <= 32'b111100_00000000000000001110000001; 	// j
disk[882] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[883] <= 32'b010000_00000_11000_0000000000000011; 	// li
disk[884] <= 32'b000000_00101_11000_10111_00000_010000; 	// gt
disk[885] <= 32'b010101_10111_00000_0000001101111010; 	// jf
disk[886] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[887] <= 32'b010010_11110_00110_1111111111111110; 	// sw
disk[888] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[889] <= 32'b111100_00000000000000001110000001; 	// j
disk[890] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[891] <= 32'b010000_00000_10000_0000000000000001; 	// li
disk[892] <= 32'b000000_00101_10000_01111_00000_001110; 	// lt
disk[893] <= 32'b010101_01111_00000_0000001110000001; 	// jf
disk[894] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[895] <= 32'b010010_11110_00110_1111111111111110; 	// sw
disk[896] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[897] <= 32'b111100_00000000000000001110111100; 	// j
disk[898] <= 32'b001111_11101_00101_0000000010101010; 	// lw
disk[899] <= 32'b001111_11101_00110_0000000010100110; 	// lw
disk[900] <= 32'b000000_00101_00110_10001_00000_001100; 	// eq
disk[901] <= 32'b010101_10001_00000_0000001110011111; 	// jf
disk[902] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[903] <= 32'b010000_00000_10011_0000000000000001; 	// li
disk[904] <= 32'b000000_00111_10011_10010_00000_001100; 	// eq
disk[905] <= 32'b010101_10010_00000_0000001110010000; 	// jf
disk[906] <= 32'b111110_00000000000000001011011101; 	// jal
disk[907] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[908] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[909] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[910] <= 32'b010010_11110_00110_1111111111111110; 	// sw
disk[911] <= 32'b111100_00000000000000001110011110; 	// j
disk[912] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[913] <= 32'b010000_00000_10101_0000000000000010; 	// li
disk[914] <= 32'b000000_00101_10101_10100_00000_001100; 	// eq
disk[915] <= 32'b010101_10100_00000_0000001110011100; 	// jf
disk[916] <= 32'b111110_00000000000000000110010100; 	// jal
disk[917] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[918] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[919] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[920] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[921] <= 32'b001111_11101_00110_0000000010101000; 	// lw
disk[922] <= 32'b010010_11110_00110_1111111111111110; 	// sw
disk[923] <= 32'b111100_00000000000000001110011110; 	// j
disk[924] <= 32'b001111_11101_00101_0000000010100011; 	// lw
disk[925] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[926] <= 32'b111100_00000000000000001110111100; 	// j
disk[927] <= 32'b001111_11101_00101_0000000010101010; 	// lw
disk[928] <= 32'b001111_11101_00110_0000000010100111; 	// lw
disk[929] <= 32'b000000_00101_00110_10110_00000_001100; 	// eq
disk[930] <= 32'b010101_10110_00000_0000001110101110; 	// jf
disk[931] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[932] <= 32'b010000_00000_11000_0000000000000000; 	// li
disk[933] <= 32'b000000_00111_11000_10111_00000_010000; 	// gt
disk[934] <= 32'b010101_10111_00000_0000001110101011; 	// jf
disk[935] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[936] <= 32'b111110_00000000000000001000110110; 	// jal
disk[937] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[938] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[939] <= 32'b001111_11101_00101_0000000010100011; 	// lw
disk[940] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[941] <= 32'b111100_00000000000000001110111100; 	// j
disk[942] <= 32'b001111_11101_00101_0000000010101010; 	// lw
disk[943] <= 32'b001111_11101_00110_0000000010101000; 	// lw
disk[944] <= 32'b000000_00101_00110_01111_00000_001100; 	// eq
disk[945] <= 32'b010101_01111_00000_0000001110111100; 	// jf
disk[946] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[947] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[948] <= 32'b000000_00111_10001_10000_00000_010000; 	// gt
disk[949] <= 32'b010101_10000_00000_0000001110111010; 	// jf
disk[950] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[951] <= 32'b111110_00000000000000001011010001; 	// jal
disk[952] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[953] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[954] <= 32'b001111_11101_00101_0000000010100011; 	// lw
disk[955] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[956] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[957] <= 32'b010010_11101_00101_0000000010101010; 	// sw
disk[958] <= 32'b001111_11101_00110_0000000010101010; 	// lw
disk[959] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[960] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[961] <= 32'b111100_00000000000000001100101001; 	// j
disk[962] <= 32'b111111_00000000000000000000000000; 	// halt


		// PROGRAMA 1
		disk[1700] <= 32'b111101_00000000000000000000100011;		// Jump to Main
		disk[1701] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[1702] <= 32'b010010_11110_00001_1111111111111100; 	// sw
		disk[1703] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[1704] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[1705] <= 32'b010000_00000_10000_0000000000000001; 	// li
		disk[1706] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[1707] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[1708] <= 32'b010010_11110_10001_1111111111111101; 	// sw
		disk[1709] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[1710] <= 32'b001111_11110_00110_1111111111111100; 	// lw
		disk[1711] <= 32'b000000_00101_00110_10010_00000_001111; 	// let
		disk[1712] <= 32'b010101_10010_00000_0000000000100000; 	// jf
		disk[1713] <= 32'b010000_00000_10100_0000000000000001; 	// li
		disk[1714] <= 32'b000000_00101_10100_10011_00000_001111; 	// let
		disk[1715] <= 32'b010101_10011_00000_0000000000010010; 	// jf
		disk[1716] <= 32'b010010_11110_00101_1111111111111110; 	// sw
		disk[1717] <= 32'b111100_00000000000000000000011011; 	// j
		disk[1718] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1719] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[1720] <= 32'b000000_00101_00110_10101_00000_000000; 	// add
		disk[1721] <= 32'b010010_11110_10101_1111111111111110; 	// sw
		disk[1722] <= 32'b010010_11110_00110_1111111111111111; 	// sw
		disk[1723] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1724] <= 32'b001111_11110_00111_1111111111111110; 	// lw
		disk[1725] <= 32'b010010_11110_00111_0000000000000000; 	// sw
		disk[1726] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[1727] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[1728] <= 32'b000001_00101_10110_0000000000000001; 	// addi
		disk[1729] <= 32'b010010_11110_10110_1111111111111101; 	// sw
		disk[1730] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[1731] <= 32'b111100_00000000000000000000001001; 	// j
		disk[1732] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[1733] <= 32'b001110_00101_11001_0000000000000000; 	// mov
		disk[1734] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1735] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[1736] <= 32'b010000_00000_01111_0000000000001011; 	// li
		disk[1737] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[1738] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1739] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1740] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1741] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[1742] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[1743] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1744] <= 32'b001110_11001_00101_0000000000000000; 	// mov
		disk[1745] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1746] <= 32'b010000_00000_00010_0000000000000000; 	// li
		disk[1747] <= 32'b010100_00000_00001_0000000000000000; 	// out
		disk[1748] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[1749] <= 32'b011111_11111_00000_0000000000000000; 	// syscall

		// PROGRAMA 2
		disk[1800] <= 32'b111101_00000000000000000000100001;		// Jump to Main
		disk[1801] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[1802] <= 32'b010010_11110_00001_1111111111111100; 	// sw
		disk[1803] <= 32'b010010_11110_00010_1111111111111101; 	// sw
		disk[1804] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[1805] <= 32'b010010_11110_01111_1111111111111110; 	// sw
		disk[1806] <= 32'b010000_00000_10000_0000000000000000; 	// li
		disk[1807] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[1808] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[1809] <= 32'b001111_11110_00110_1111111111111101; 	// lw
		disk[1810] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
		disk[1811] <= 32'b010101_10001_00000_0000000000011100; 	// jf
		disk[1812] <= 32'b001111_11110_00111_1111111111111100; 	// lw
		disk[1813] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
		disk[1814] <= 32'b001111_10010_10010_0000000000000000; 	// lw
		disk[1815] <= 32'b001111_11110_01000_0000000000000000; 	// lw
		disk[1816] <= 32'b000000_01000_10010_10011_00000_001110; 	// lt
		disk[1817] <= 32'b010101_10011_00000_0000000000010111; 	// jf
		disk[1818] <= 32'b000000_00111_00101_10100_00000_000000; 	// add
		disk[1819] <= 32'b001111_10100_10100_0000000000000000; 	// lw
		disk[1820] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[1821] <= 32'b001111_11110_01000_0000000000000000; 	// lw
		disk[1822] <= 32'b010010_11110_00101_1111111111111111; 	// sw
		disk[1823] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[1824] <= 32'b000001_00101_10101_0000000000000001; 	// addi
		disk[1825] <= 32'b010010_11110_10101_1111111111111110; 	// sw
		disk[1826] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[1827] <= 32'b111100_00000000000000000000001000; 	// j
		disk[1828] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1829] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1830] <= 32'b010000_00000_00010_0000000000000001; 	// li
		disk[1831] <= 32'b010100_00000_00001_0000000000000001; 	// out
		disk[1832] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1833] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[1834] <= 32'b010001_11110_00101_1111111111111011; 	// la
		disk[1835] <= 32'b010000_00000_01111_0000000000001100; 	// li
		disk[1836] <= 32'b010010_00101_01111_0000000000000000; 	// sw
		disk[1837] <= 32'b010000_00000_10000_0000000000101001; 	// li
		disk[1838] <= 32'b010010_00101_10000_0000000000000001; 	// sw
		disk[1839] <= 32'b010000_00000_10001_0000000000010111; 	// li
		disk[1840] <= 32'b010010_00101_10001_0000000000000010; 	// sw
		disk[1841] <= 32'b010000_00000_10010_0000000001100010; 	// li
		disk[1842] <= 32'b010010_00101_10010_0000000000000011; 	// sw
		disk[1843] <= 32'b010000_00000_10011_0000000000100001; 	// li
		disk[1844] <= 32'b010010_00101_10011_0000000000000100; 	// sw
		disk[1845] <= 32'b010000_00000_10100_0000000000010101; 	// li
		disk[1846] <= 32'b010010_00101_10100_0000000000000101; 	// sw
		disk[1847] <= 32'b010001_11110_00001_1111111111111011; 	// la
		disk[1848] <= 32'b010000_00000_00010_0000000000000110; 	// li
		disk[1849] <= 32'b010010_11110_11111_1111111111111010; 	// sw
		disk[1850] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[1851] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[1852] <= 32'b001111_11110_11111_1111111111111010; 	// lw
		disk[1853] <= 32'b001110_11001_00101_0000000000000000; 	// mov
		disk[1854] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[1855] <= 32'b011111_11111_00000_0000000000000000; 	// syscall
		
		// PROGRAMA 3
		disk[1900] <= 32'b111101_00000000000000000000010100;		// Jump to Main
		disk[1901] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[1902] <= 32'b010010_11110_00001_1111111111111111; 	// sw
		disk[1903] <= 32'b010000_00000_01111_0000000000000001; 	// li
		disk[1904] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[1905] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1906] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[1907] <= 32'b000000_00101_10001_10000_00000_010000; 	// gt
		disk[1908] <= 32'b010101_10000_00000_0000000000010001; 	// jf
		disk[1909] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[1910] <= 32'b000000_00110_00101_10010_00000_000010; 	// mul
		disk[1911] <= 32'b010010_11110_10010_0000000000000000; 	// sw
		disk[1912] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[1913] <= 32'b000010_00101_10011_0000000000000001; 	// subi
		disk[1914] <= 32'b010010_11110_10011_1111111111111111; 	// sw
		disk[1915] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1916] <= 32'b111100_00000000000000000000000101; 	// j
		disk[1917] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1918] <= 32'b001110_00101_11001_0000000000000000; 	// mov
		disk[1919] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1920] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[1921] <= 32'b101000_00000000000000000000000000; 	// preIO
		disk[1922] <= 32'b010011_00000_01111_0000000000000000; 	// in
		disk[1923] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[1924] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1925] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1926] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1927] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[1928] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[1929] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1930] <= 32'b001110_11001_00101_0000000000000000; 	// mov
		disk[1931] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1932] <= 32'b010000_00000_00010_0000000000000010; 	// li
		disk[1933] <= 32'b010100_00000_00001_0000000000000010; 	// out
		disk[1934] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[1935] <= 32'b011111_11111_00000_0000000000000000; 	// syscall

	end
endmodule
