library verilog;
use verilog.vl_types.all;
entity multiplexador_escrita_br_vlg_vec_tst is
end multiplexador_escrita_br_vlg_vec_tst;
