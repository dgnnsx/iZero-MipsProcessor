module disco_rigido(pc, instrucao);
	// Entrada
	input [25:0] pc;				// PC Atual
	
	// Saida
	output [31:0] instrucao;	// Proxima instrucao a ser executada
	
	parameter DISK_SIZE = 71; // Tamanho do disco
	wire [31:0] disk [DISK_SIZE-1:0];

	assign disk[0] = 32'b010110_00000000000000000000100001;		// Jump to Main
	assign disk[1] = 32'b000001_11110_11110_0000000000000011; 	// addi
	assign disk[2] = 32'b010010_11110_00110_0000000000000000; 	// sw
	assign disk[3] = 32'b001111_11110_01010_0000000000000000; 	// lw
	assign disk[4] = 32'b010000_00000_10101_0000000000000010; 	// li
	assign disk[5] = 32'b000000_01010_10101_10100_00000_001110; 	// lt
	assign disk[6] = 32'b010101_10100_00000_0000000000001010; 	// jf
	assign disk[7] = 32'b010000_00000_10110_0000000000000001; 	// li
	assign disk[8] = 32'b001110_10110_00001_0000000000000000; 	// mov
	assign disk[9] = 32'b000000_11111_00000_00000_00000_010010; 	// jr
	assign disk[10] = 32'b000010_01010_10111_0000000000000001; 	// subi
	assign disk[11] = 32'b001110_10111_00110_0000000000000000; 	// mov
	assign disk[12] = 32'b010010_11110_11111_1111111111111110; 	// sw
	assign disk[13] = 32'b010010_11110_01010_0000000000000000; 	// sw
	assign disk[14] = 32'b010111_00000000000000000000000001; 	// jal
	assign disk[15] = 32'b000010_11110_11110_0000000000000011; 	// subi
	assign disk[16] = 32'b001111_11110_11111_1111111111111110; 	// lw
	assign disk[17] = 32'b001111_11110_01010_0000000000000000; 	// lw
	assign disk[18] = 32'b001110_00001_01011_0000000000000000; 	// mov
	assign disk[19] = 32'b000010_01010_11000_0000000000000010; 	// subi
	assign disk[20] = 32'b001110_11000_00110_0000000000000000; 	// mov
	assign disk[21] = 32'b010010_11110_11111_1111111111111110; 	// sw
	assign disk[22] = 32'b010010_11110_01010_0000000000000000; 	// sw
	assign disk[23] = 32'b010010_11110_01011_1111111111111111; 	// sw
	assign disk[24] = 32'b010111_00000000000000000000000001; 	// jal
	assign disk[25] = 32'b000010_11110_11110_0000000000000011; 	// subi
	assign disk[26] = 32'b001111_11110_11111_1111111111111110; 	// lw
	assign disk[27] = 32'b001111_11110_01010_0000000000000000; 	// lw
	assign disk[28] = 32'b001111_11110_01011_1111111111111111; 	// lw
	assign disk[29] = 32'b001110_00001_01100_0000000000000000; 	// mov
	assign disk[30] = 32'b000000_01011_01100_11001_00000_000000; 	// add
	assign disk[31] = 32'b001110_11001_00001_0000000000000000; 	// mov
	assign disk[32] = 32'b000000_11111_00000_00000_00000_010010; 	// jr
	assign disk[33] = 32'b000001_11110_11110_0000000000000001; 	// addi
	assign disk[34] = 32'b010011_00000_10100_0000000000000000; 	// in
	assign disk[35] = 32'b010010_11110_10100_0000000000000000; 	// sw
	assign disk[36] = 32'b001111_11110_01010_0000000000000000; 	// lw
	assign disk[37] = 32'b001110_01010_00110_0000000000000000; 	// mov
	assign disk[38] = 32'b010010_11110_01010_0000000000000000; 	// sw
	assign disk[39] = 32'b010111_00000000000000000000000001; 	// jal
	assign disk[40] = 32'b001110_00001_01011_0000000000000000; 	// mov
	assign disk[41] = 32'b000010_11110_11110_0000000000000011; 	// subi
	assign disk[42] = 32'b001111_11110_01010_0000000000000000; 	// lw
	assign disk[43] = 32'b001110_01011_00110_0000000000000000; 	// mov
	assign disk[44] = 32'b010000_00000_00111_0000000000000010; 	// li
	assign disk[45] = 32'b010100_00000_00110_0000000000000010; 	// out
	assign disk[46] = 32'b011000_00000000000000000000000000; 	// halt

	assign instrucao = pc < DISK_SIZE ? disk[pc] : disk[DISK_SIZE-1];
endmodule
