library verilog;
use verilog.vl_types.all;
entity unidade_logica_aritmetica_vlg_vec_tst is
end unidade_logica_aritmetica_vlg_vec_tst;
