module memoria_de_instrucoes(pc, instrucao);
	// Entrada
	input [25:0] pc;				// PC Atual
	
	// Saida
	output [31:0] instrucao;	// Proxima instrucao a ser executada
	
	parameter MEM_SIZE = 150; // Tamanho da memoria
	wire [31:0] rom [MEM_SIZE-1:0];// Memoria de instrucoes

	assign rom[0] = 32'b010110_00000000000000000000100110;		// Jump to Main
assign rom[1] = 32'b000001_11110_11110_0000000000000100; 	// addi
assign rom[2] = 32'b010010_11110_00110_1111111111111110; 	// sw
assign rom[3] = 32'b001111_11110_01010_1111111111111110; 	// lw
assign rom[4] = 32'b010000_00000_10101_0000000000000000; 	// li
assign rom[5] = 32'b000000_01010_10101_10100_00000_001100; 	// lt
assign rom[6] = 32'b010101_10100_00000_0000000000001010; 	// jf
assign rom[7] = 32'b010000_00000_10110_0000000000000000; 	// li
assign rom[8] = 32'b001110_10110_00001_0000000000000000; 	// mov
assign rom[9] = 32'b000000_11111_00000_00000_00000_010010; 	// jr
assign rom[10] = 32'b010000_00000_11000_0000000000000001; 	// li
assign rom[11] = 32'b000000_01010_11000_10111_00000_001100; 	// lt
assign rom[12] = 32'b010101_10111_00000_0000000000010000; 	// jf
assign rom[13] = 32'b010000_00000_11001_0000000000000001; 	// li
assign rom[14] = 32'b001110_11001_00001_0000000000000000; 	// mov
assign rom[15] = 32'b000000_11111_00000_00000_00000_010010; 	// jr
assign rom[16] = 32'b000010_01010_11010_0000000000000001; 	// subi
assign rom[17] = 32'b001110_11010_00110_0000000000000000; 	// mov
assign rom[18] = 32'b010010_11110_11111_0000000000000001; 	// sw
assign rom[19] = 32'b010111_00000000000000000000000001; 	// jal
assign rom[20] = 32'b000010_11110_11110_0000000000000100; 	// subi
assign rom[21] = 32'b001111_11110_11111_0000000000000001; 	// lw
assign rom[22] = 32'b001110_00001_11011_0000000000000000; 	// mov
assign rom[23] = 32'b010010_11110_11011_1111111111111111; 	// sw
assign rom[24] = 32'b001111_11110_01010_1111111111111110; 	// lw
assign rom[25] = 32'b000010_01010_11100_0000000000000010; 	// subi
assign rom[26] = 32'b001110_11100_00110_0000000000000000; 	// mov
assign rom[27] = 32'b010010_11110_11111_0000000000000001; 	// sw
assign rom[28] = 32'b010111_00000000000000000000000001; 	// jal
assign rom[29] = 32'b000010_11110_11110_0000000000000100; 	// subi
assign rom[30] = 32'b001111_11110_11111_0000000000000001; 	// lw
assign rom[31] = 32'b001110_00001_11101_0000000000000000; 	// mov
assign rom[32] = 32'b010010_11110_11101_0000000000000000; 	// sw
assign rom[33] = 32'b001111_11110_01010_1111111111111111; 	// lw
assign rom[34] = 32'b001111_11110_01011_0000000000000000; 	// lw
assign rom[35] = 32'b000000_01010_01011_10100_00000_000000; 	// add
assign rom[36] = 32'b001110_10100_00001_0000000000000000; 	// mov
assign rom[37] = 32'b000000_11111_00000_00000_00000_010010; 	// jr
assign rom[38] = 32'b000001_11110_11110_0000000000000001; 	// addi
assign rom[39] = 32'b010011_00000_10100_0000000000000000; 	// in
assign rom[40] = 32'b010010_11110_10100_0000000000000000; 	// sw
assign rom[41] = 32'b001111_11110_01010_0000000000000000; 	// lw
assign rom[42] = 32'b001110_01010_00110_0000000000000000; 	// mov
assign rom[43] = 32'b010111_00000000000000000000000001; 	// jal
assign rom[44] = 32'b001110_00001_10101_0000000000000000; 	// mov
assign rom[45] = 32'b000010_11110_11110_0000000000000100; 	// subi
assign rom[46] = 32'b001110_10101_00110_0000000000000000; 	// mov
assign rom[47] = 32'b010000_00000_00111_0000000000000010; 	// li
assign rom[48] = 32'b010100_00000_00110_0000000000000010; 	// out
assign rom[49] = 32'b011000_00000000000000000000000000; 	// halt
	assign instrucao = rom[pc];
endmodule
