library verilog;
use verilog.vl_types.all;
entity BCD_quatro_digitos_vlg_vec_tst is
end BCD_quatro_digitos_vlg_vec_tst;
