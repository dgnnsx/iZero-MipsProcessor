module disco_rigido (clk, we, addr, datain, dataout);
	input clk;										// clock
	input we;										// write enable
	input [31:0] addr;							// disk address
	input [31:0] datain;							// data in (to disk)
	
	output reg [31:0] dataout;					// data out (from disk)
	
	localparam DISK_SIZE = 4096;				// Tamanho do disco
	reg [31:0] disk [DISK_SIZE-1:0];			// disk cells
	
	always @ (posedge clk) begin
		if (we) disk[addr] <= datain;			// write disk
	end
	
	always @ (negedge clk) begin
		dataout <= disk[addr];
	end

	initial begin
		// SISTEMA OPERACIONAL

disk[0] <= 32'b111100_00000000000000010101110110;		// Jump to Main
disk[1] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[2] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[3] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[4] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[5] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[6] <= 32'b010110_00001_10000_0000000000000000; 	// ldk
disk[7] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[8] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[9] <= 32'b001101_00101_10001_0000000000011010; 	// srli
disk[10] <= 32'b001111_11101_00110_0000000110101010; 	// lw
disk[11] <= 32'b000000_10001_00110_10010_00000_001101; 	// ne
disk[12] <= 32'b010101_10010_00000_0000000000010110; 	// jf
disk[13] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[14] <= 32'b000001_00111_10011_0000000000000001; 	// addi
disk[15] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[16] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[17] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[18] <= 32'b010110_00001_10100_0000000000000000; 	// ldk
disk[19] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[20] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[21] <= 32'b111100_00000000000000000000001000; 	// j
disk[22] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[23] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[24] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[25] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[26] <= 32'b010010_11110_00001_1111111111111111; 	// sw
disk[27] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[28] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[29] <= 32'b000000_00101_10000_01111_00000_001100; 	// eq
disk[30] <= 32'b010101_01111_00000_0000000000100010; 	// jf
disk[31] <= 32'b010000_00000_10001_0000000000000001; 	// li
disk[32] <= 32'b001110_10001_11000_0000000000000000; 	// mov
disk[33] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[34] <= 32'b010000_00000_10010_0000000000000001; 	// li
disk[35] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[36] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[37] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[38] <= 32'b000000_00101_10100_10011_00000_010000; 	// gt
disk[39] <= 32'b010101_10011_00000_0000000000110000; 	// jf
disk[40] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[41] <= 32'b000011_00110_10101_0000000000000010; 	// muli
disk[42] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[43] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[44] <= 32'b000010_00101_10110_0000000000000001; 	// subi
disk[45] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[46] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[47] <= 32'b111100_00000000000000000000100100; 	// j
disk[48] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[49] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[50] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[51] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[52] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[53] <= 32'b010000_00000_00010_0000000000000000; 	// li
disk[54] <= 32'b010100_00000_00001_0000000000000000; 	// out
disk[55] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[56] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[57] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[58] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[59] <= 32'b010000_00000_00010_0000000000000010; 	// li
disk[60] <= 32'b010100_00000_00001_0000000000000010; 	// out
disk[61] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[62] <= 32'b000001_11110_11110_0000000000000110; 	// addi
disk[63] <= 32'b010001_11101_00101_0000000001000000; 	// la
disk[64] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[65] <= 32'b000000_00101_00110_01111_00000_000000; 	// add
disk[66] <= 32'b001111_01111_01111_0000000000000000; 	// lw
disk[67] <= 32'b000001_01111_10000_0000000000000001; 	// addi
disk[68] <= 32'b010010_11110_10000_1111111111111110; 	// sw
disk[69] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[70] <= 32'b001111_11101_01000_0000000011101011; 	// lw
disk[71] <= 32'b000000_00111_01000_10001_00000_000010; 	// mul
disk[72] <= 32'b010010_11110_10001_1111111111111111; 	// sw
disk[73] <= 32'b001111_11101_01001_0000000011101100; 	// lw
disk[74] <= 32'b000010_01001_10010_0000000000000001; 	// subi
disk[75] <= 32'b000000_01000_10010_10011_00000_000010; 	// mul
disk[76] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[77] <= 32'b001111_11101_00101_0000000011101011; 	// lw
disk[78] <= 32'b001111_11101_00110_0000000011101100; 	// lw
disk[79] <= 32'b000000_00101_00110_10100_00000_000010; 	// mul
disk[80] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[81] <= 32'b000000_00111_10100_10101_00000_001110; 	// lt
disk[82] <= 32'b010101_10101_00000_0000000001100010; 	// jf
disk[83] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[84] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[85] <= 32'b001111_00001_10110_0000000000000000; 	// lw
disk[86] <= 32'b010010_11110_10110_1111111111111101; 	// sw
disk[87] <= 32'b001111_11110_01001_1111111111111101; 	// lw
disk[88] <= 32'b001110_01001_00001_0000000000000000; 	// mov
disk[89] <= 32'b001110_00111_00010_0000000000000000; 	// mov
disk[90] <= 32'b010010_00010_00001_0000000000000000; 	// sw
disk[91] <= 32'b000001_01000_10111_0000000000000001; 	// addi
disk[92] <= 32'b010010_11110_10111_1111111111111111; 	// sw
disk[93] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[94] <= 32'b000001_00111_01111_0000000000000001; 	// addi
disk[95] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[96] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[97] <= 32'b111100_00000000000000000001001101; 	// j
disk[98] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[99] <= 32'b000001_11110_11110_0000000000000110; 	// addi
disk[100] <= 32'b010010_11110_00001_1111111111111101; 	// sw
disk[101] <= 32'b001111_11110_00101_1111111111111101; 	// lw
disk[102] <= 32'b000001_00101_01111_0000000000000001; 	// addi
disk[103] <= 32'b010010_11110_01111_1111111111111101; 	// sw
disk[104] <= 32'b001111_11110_00101_1111111111111101; 	// lw
disk[105] <= 32'b001111_11101_00110_0000000011101100; 	// lw
disk[106] <= 32'b000010_00110_10000_0000000000000001; 	// subi
disk[107] <= 32'b001111_11101_00111_0000000011101011; 	// lw
disk[108] <= 32'b000000_00111_10000_10001_00000_000010; 	// mul
disk[109] <= 32'b010010_11110_10001_1111111111111111; 	// sw
disk[110] <= 32'b000000_00101_00111_10010_00000_000010; 	// mul
disk[111] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[112] <= 32'b001111_11101_00101_0000000011101011; 	// lw
disk[113] <= 32'b001111_11101_00110_0000000011101100; 	// lw
disk[114] <= 32'b000000_00101_00110_10011_00000_000010; 	// mul
disk[115] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[116] <= 32'b000000_00111_10011_10100_00000_001110; 	// lt
disk[117] <= 32'b010101_10100_00000_0000000010000101; 	// jf
disk[118] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[119] <= 32'b001111_00001_10101_0000000000000000; 	// lw
disk[120] <= 32'b010010_11110_10101_1111111111111110; 	// sw
disk[121] <= 32'b001111_11110_01000_1111111111111110; 	// lw
disk[122] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[123] <= 32'b001111_11110_01001_0000000000000000; 	// lw
disk[124] <= 32'b001110_01001_00010_0000000000000000; 	// mov
disk[125] <= 32'b010010_00010_00001_0000000000000000; 	// sw
disk[126] <= 32'b000001_00111_10110_0000000000000001; 	// addi
disk[127] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[128] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[129] <= 32'b000001_01001_10111_0000000000000001; 	// addi
disk[130] <= 32'b010010_11110_10111_0000000000000000; 	// sw
disk[131] <= 32'b001111_11110_01001_0000000000000000; 	// lw
disk[132] <= 32'b111100_00000000000000000001110000; 	// j
disk[133] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[134] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[135] <= 32'b010010_11110_00001_1111111111111110; 	// sw
disk[136] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[137] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[138] <= 32'b010010_11101_01111_0000000001011111; 	// sw
disk[139] <= 32'b010001_11101_00110_0000000000110110; 	// la
disk[140] <= 32'b001111_11101_00111_0000000001011111; 	// lw
disk[141] <= 32'b000000_00110_00111_10000_00000_000000; 	// add
disk[142] <= 32'b001111_10000_10000_0000000000000000; 	// lw
disk[143] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[144] <= 32'b010001_11101_01000_0000000001001010; 	// la
disk[145] <= 32'b000000_01000_00111_10001_00000_000000; 	// add
disk[146] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[147] <= 32'b010010_11110_10001_0000000000000000; 	// sw
disk[148] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[149] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[150] <= 32'b000000_00101_10011_10010_00000_010000; 	// gt
disk[151] <= 32'b010101_10010_00000_0000000010100100; 	// jf
disk[152] <= 32'b010001_11101_00110_0000000001101011; 	// la
disk[153] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[154] <= 32'b000000_00110_00111_10100_00000_000000; 	// add
disk[155] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[156] <= 32'b010010_10100_10101_0000000000000000; 	// sw
disk[157] <= 32'b000001_00111_10110_0000000000000001; 	// addi
disk[158] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[159] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[160] <= 32'b000010_00101_10111_0000000000000001; 	// subi
disk[161] <= 32'b010010_11110_10111_0000000000000000; 	// sw
disk[162] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[163] <= 32'b111100_00000000000000000010010100; 	// j
disk[164] <= 32'b010001_11101_00101_0000000110010100; 	// la
disk[165] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[166] <= 32'b000000_00101_00110_01111_00000_000000; 	// add
disk[167] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[168] <= 32'b010010_01111_10000_0000000000000000; 	// sw
disk[169] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[170] <= 32'b000000_00111_00110_10001_00000_000000; 	// add
disk[171] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[172] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[173] <= 32'b010001_11101_01000_0000000000001110; 	// la
disk[174] <= 32'b000000_01000_00110_10011_00000_000000; 	// add
disk[175] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[176] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[177] <= 32'b010001_11101_01001_0000000000011000; 	// la
disk[178] <= 32'b000000_01001_00110_10101_00000_000000; 	// add
disk[179] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[180] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[181] <= 32'b010001_11101_01010_0000000000100010; 	// la
disk[182] <= 32'b000000_01010_00110_10111_00000_000000; 	// add
disk[183] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[184] <= 32'b010010_10111_01111_0000000000000000; 	// sw
disk[185] <= 32'b010001_11101_01011_0000000000101100; 	// la
disk[186] <= 32'b000000_01011_00110_10000_00000_000000; 	// add
disk[187] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[188] <= 32'b010010_10000_10001_0000000000000000; 	// sw
disk[189] <= 32'b010001_11101_01100_0000000001000000; 	// la
disk[190] <= 32'b000000_01100_00110_10010_00000_000000; 	// add
disk[191] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[192] <= 32'b010010_10010_10011_0000000000000000; 	// sw
disk[193] <= 32'b010001_11101_01101_0000000001001010; 	// la
disk[194] <= 32'b000000_01101_00110_10100_00000_000000; 	// add
disk[195] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[196] <= 32'b010010_10100_10101_0000000000000000; 	// sw
disk[197] <= 32'b010001_11101_01110_0000000001010100; 	// la
disk[198] <= 32'b000000_01110_00110_10110_00000_000000; 	// add
disk[199] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[200] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[201] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[202] <= 32'b010010_11101_01111_0000000001011111; 	// sw
disk[203] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[204] <= 32'b010000_00000_10000_0000001111100111; 	// li
disk[205] <= 32'b010010_11101_10000_0000000001011110; 	// sw
disk[206] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[207] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[208] <= 32'b010010_11110_00001_1111111111111110; 	// sw
disk[209] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[210] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[211] <= 32'b010010_11110_01111_1111111111111110; 	// sw
disk[212] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[213] <= 32'b010001_11101_00110_0000000000000100; 	// la
disk[214] <= 32'b000000_00110_00101_10000_00000_000000; 	// add
disk[215] <= 32'b001111_10000_10000_0000000000000000; 	// lw
disk[216] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[217] <= 32'b000000_10000_10010_10001_00000_001101; 	// ne
disk[218] <= 32'b010101_10001_00000_0000000011100010; 	// jf
disk[219] <= 32'b000001_00101_10011_0000000000000001; 	// addi
disk[220] <= 32'b001110_10011_00001_0000000000000000; 	// mov
disk[221] <= 32'b010010_11110_11111_1111111111111101; 	// sw
disk[222] <= 32'b111110_00000000000000000010000110; 	// jal
disk[223] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[224] <= 32'b001111_11110_11111_1111111111111101; 	// lw
disk[225] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[226] <= 32'b010001_11101_00101_0000000110000000; 	// la
disk[227] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[228] <= 32'b000000_00101_00110_10100_00000_000000; 	// add
disk[229] <= 32'b001111_10100_10100_0000000000000000; 	// lw
disk[230] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[231] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[232] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[233] <= 32'b010110_00001_10101_0000000000000000; 	// ldk
disk[234] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[235] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[236] <= 32'b001101_00101_10110_0000000000011010; 	// srli
disk[237] <= 32'b001111_11101_00110_0000000110101000; 	// lw
disk[238] <= 32'b000000_10110_00110_10111_00000_001101; 	// ne
disk[239] <= 32'b010101_10111_00000_0000000011111100; 	// jf
disk[240] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[241] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[242] <= 32'b001110_00111_00010_0000000000000000; 	// mov
disk[243] <= 32'b010111_00010_00001_0000000000000000; 	// sdk
disk[244] <= 32'b000001_00111_01111_0000000000000001; 	// addi
disk[245] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[246] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[247] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[248] <= 32'b010110_00001_10000_0000000000000000; 	// ldk
disk[249] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[250] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[251] <= 32'b111100_00000000000000000011101011; 	// j
disk[252] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[253] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[254] <= 32'b001110_00101_00010_0000000000000000; 	// mov
disk[255] <= 32'b010111_00010_00001_0000000000000000; 	// sdk
disk[256] <= 32'b010001_11101_00110_0000000101110110; 	// la
disk[257] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[258] <= 32'b000000_00110_00111_10001_00000_000000; 	// add
disk[259] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[260] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[261] <= 32'b010001_11101_01000_0000000110001010; 	// la
disk[262] <= 32'b000000_01000_00111_10011_00000_000000; 	// add
disk[263] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[264] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[265] <= 32'b010001_11101_01001_0000000110000000; 	// la
disk[266] <= 32'b000000_01001_00111_10101_00000_000000; 	// add
disk[267] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[268] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[269] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[270] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[271] <= 32'b010010_11110_00001_1111111111111111; 	// sw
disk[272] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[273] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[274] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[275] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[276] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[277] <= 32'b100100_00000_00001_0000000000000000; 	// lcdCurr
disk[278] <= 32'b001111_11101_00110_0000000110110101; 	// lw
disk[279] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[280] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[281] <= 32'b010011_00000_10000_0000000000000000; 	// in
disk[282] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[283] <= 32'b010001_11101_00111_0000000110001010; 	// la
disk[284] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[285] <= 32'b001111_11110_01000_0000000000000000; 	// lw
disk[286] <= 32'b010010_10001_01000_0000000000000000; 	// sw
disk[287] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[288] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[289] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[290] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[291] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[292] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[293] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[294] <= 32'b001111_11101_00110_0000000011101110; 	// lw
disk[295] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[296] <= 32'b010101_10001_00000_0000000101000010; 	// jf
disk[297] <= 32'b010001_11101_00111_0000000101110110; 	// la
disk[298] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
disk[299] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[300] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[301] <= 32'b000000_10010_10100_10011_00000_001101; 	// ne
disk[302] <= 32'b010101_10011_00000_0000000100111101; 	// jf
disk[303] <= 32'b010001_11101_01000_0000000110001010; 	// la
disk[304] <= 32'b000000_01000_00101_10101_00000_000000; 	// add
disk[305] <= 32'b001111_10101_10101_0000000000000000; 	// lw
disk[306] <= 32'b000010_10101_10110_0000000000000001; 	// subi
disk[307] <= 32'b001110_10110_00001_0000000000000000; 	// mov
disk[308] <= 32'b010010_11110_11111_1111111111111110; 	// sw
disk[309] <= 32'b111110_00000000000000000000011001; 	// jal
disk[310] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[311] <= 32'b001111_11110_11111_1111111111111110; 	// lw
disk[312] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[313] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[314] <= 32'b000000_00110_00101_10111_00000_000000; 	// add
disk[315] <= 32'b010010_11110_10111_0000000000000000; 	// sw
disk[316] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[317] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[318] <= 32'b000001_00101_01111_0000000000000001; 	// addi
disk[319] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[320] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[321] <= 32'b111100_00000000000000000100100101; 	// j
disk[322] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[323] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[324] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[325] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[326] <= 32'b010000_00000_01111_0000000000000010; 	// li
disk[327] <= 32'b010010_11101_01111_0000000101110100; 	// sw
disk[328] <= 32'b010000_00000_10000_0000000000000001; 	// li
disk[329] <= 32'b010010_11101_10000_0000000101110101; 	// sw
disk[330] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[331] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[332] <= 32'b010000_00000_01111_0000000000000001; 	// li
disk[333] <= 32'b010010_11101_01111_0000000000000000; 	// sw
disk[334] <= 32'b010000_00000_10000_0000000000000010; 	// li
disk[335] <= 32'b010010_11101_10000_0000000000000001; 	// sw
disk[336] <= 32'b010000_00000_10001_0000000000000011; 	// li
disk[337] <= 32'b010010_11101_10001_0000000000000010; 	// sw
disk[338] <= 32'b010000_00000_10010_0000000110010100; 	// li
disk[339] <= 32'b010010_11101_10010_0000000000000011; 	// sw
disk[340] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[341] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[342] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[343] <= 32'b010000_00000_10101_0000000000001010; 	// li
disk[344] <= 32'b000000_00101_10101_10100_00000_001110; 	// lt
disk[345] <= 32'b010101_10100_00000_0000000110000010; 	// jf
disk[346] <= 32'b010001_11101_00110_0000000000000100; 	// la
disk[347] <= 32'b000000_00110_00101_10110_00000_000000; 	// add
disk[348] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[349] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[350] <= 32'b010001_11101_00111_0000000000001110; 	// la
disk[351] <= 32'b000000_00111_00101_01111_00000_000000; 	// add
disk[352] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[353] <= 32'b010010_01111_10000_0000000000000000; 	// sw
disk[354] <= 32'b010001_11101_01000_0000000000011000; 	// la
disk[355] <= 32'b000000_01000_00101_10001_00000_000000; 	// add
disk[356] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[357] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[358] <= 32'b010001_11101_01001_0000000000100010; 	// la
disk[359] <= 32'b000000_01001_00101_10011_00000_000000; 	// add
disk[360] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[361] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[362] <= 32'b010001_11101_01010_0000000000101100; 	// la
disk[363] <= 32'b000000_01010_00101_10101_00000_000000; 	// add
disk[364] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[365] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[366] <= 32'b010001_11101_01011_0000000001000000; 	// la
disk[367] <= 32'b000000_01011_00101_10111_00000_000000; 	// add
disk[368] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[369] <= 32'b010010_10111_01111_0000000000000000; 	// sw
disk[370] <= 32'b010001_11101_01100_0000000001001010; 	// la
disk[371] <= 32'b000000_01100_00101_10000_00000_000000; 	// add
disk[372] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[373] <= 32'b010010_10000_10001_0000000000000000; 	// sw
disk[374] <= 32'b010001_11101_01101_0000000001010100; 	// la
disk[375] <= 32'b000000_01101_00101_10010_00000_000000; 	// add
disk[376] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[377] <= 32'b010010_10010_10011_0000000000000000; 	// sw
disk[378] <= 32'b010001_11101_01110_0000000001100000; 	// la
disk[379] <= 32'b000000_01110_00101_10100_00000_000000; 	// add
disk[380] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[381] <= 32'b010010_10100_10101_0000000000000000; 	// sw
disk[382] <= 32'b000001_00101_10110_0000000000000001; 	// addi
disk[383] <= 32'b010010_11110_10110_0000000000000000; 	// sw
disk[384] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[385] <= 32'b111100_00000000000000000101010110; 	// j
disk[386] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[387] <= 32'b010010_11101_10111_0000000001101010; 	// sw
disk[388] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[389] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[390] <= 32'b010000_00000_01111_0000000000100000; 	// li
disk[391] <= 32'b010010_11101_01111_0000000011101011; 	// sw
disk[392] <= 32'b010000_00000_10000_0000000010000000; 	// li
disk[393] <= 32'b010010_11101_10000_0000000011101100; 	// sw
disk[394] <= 32'b010000_00000_10001_0000000001100100; 	// li
disk[395] <= 32'b010010_11101_10001_0000000011101101; 	// sw
disk[396] <= 32'b010000_00000_10010_0000000000001010; 	// li
disk[397] <= 32'b010010_11101_10010_0000000011101110; 	// sw
disk[398] <= 32'b010000_00000_10011_0000001111100111; 	// li
disk[399] <= 32'b010010_11101_10011_0000000001011110; 	// sw
disk[400] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[401] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[402] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[403] <= 32'b010010_11101_01111_0000000110101011; 	// sw
disk[404] <= 32'b010000_00000_10000_0000000000000001; 	// li
disk[405] <= 32'b010010_11101_10000_0000000110101100; 	// sw
disk[406] <= 32'b010000_00000_10001_0000000000000010; 	// li
disk[407] <= 32'b010010_11101_10001_0000000110101101; 	// sw
disk[408] <= 32'b010000_00000_10010_0000000000000011; 	// li
disk[409] <= 32'b010010_11101_10010_0000000110101110; 	// sw
disk[410] <= 32'b010000_00000_10011_0000000000000100; 	// li
disk[411] <= 32'b010010_11101_10011_0000000110101111; 	// sw
disk[412] <= 32'b010000_00000_10100_0000000000000101; 	// li
disk[413] <= 32'b010010_11101_10100_0000000110110000; 	// sw
disk[414] <= 32'b010000_00000_10101_0000000000000110; 	// li
disk[415] <= 32'b010010_11101_10101_0000000110110001; 	// sw
disk[416] <= 32'b010000_00000_10110_0000000000000111; 	// li
disk[417] <= 32'b010010_11101_10110_0000000110110010; 	// sw
disk[418] <= 32'b010000_00000_10111_0000000000001000; 	// li
disk[419] <= 32'b010010_11101_10111_0000000110110011; 	// sw
disk[420] <= 32'b010000_00000_01111_0000000000001001; 	// li
disk[421] <= 32'b010010_11101_01111_0000000110110100; 	// sw
disk[422] <= 32'b010000_00000_10000_0000000000011110; 	// li
disk[423] <= 32'b010010_11101_10000_0000000110110101; 	// sw
disk[424] <= 32'b001111_11101_00101_0000000110101011; 	// lw
disk[425] <= 32'b010010_11101_00101_0000000110110110; 	// sw
disk[426] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[427] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[428] <= 32'b010000_00000_01111_0000111111111111; 	// li
disk[429] <= 32'b010010_11101_01111_0000000011110000; 	// sw
disk[430] <= 32'b010000_00000_10000_0000000000011111; 	// li
disk[431] <= 32'b010010_11101_10000_0000000110101000; 	// sw
disk[432] <= 32'b010000_00000_10001_0000000000111101; 	// li
disk[433] <= 32'b010010_11101_10001_0000000110101001; 	// sw
disk[434] <= 32'b010000_00000_10010_0000000000111111; 	// li
disk[435] <= 32'b010010_11101_10010_0000000110101010; 	// sw
disk[436] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[437] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[438] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[439] <= 32'b010010_11110_01111_1111111111111110; 	// sw
disk[440] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[441] <= 32'b001111_11101_00110_0000000011101100; 	// lw
disk[442] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[443] <= 32'b010101_10000_00000_0000000111001000; 	// jf
disk[444] <= 32'b010001_11101_00111_0000000001101011; 	// la
disk[445] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[446] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[447] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[448] <= 32'b010001_11101_01000_0000000011110100; 	// la
disk[449] <= 32'b000000_01000_00101_10011_00000_000000; 	// add
disk[450] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[451] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[452] <= 32'b000001_00101_10101_0000000000000001; 	// addi
disk[453] <= 32'b010010_11110_10101_1111111111111110; 	// sw
disk[454] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[455] <= 32'b111100_00000000000000000110111000; 	// j
disk[456] <= 32'b010010_11110_11111_1111111111111101; 	// sw
disk[457] <= 32'b111110_00000000000000000000000001; 	// jal
disk[458] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[459] <= 32'b001111_11110_11111_1111111111111101; 	// lw
disk[460] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[461] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[462] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[463] <= 32'b000001_00110_10110_0000000000000001; 	// addi
disk[464] <= 32'b010010_11101_10110_0000000011101111; 	// sw
disk[465] <= 32'b001111_11101_00111_0000000011101011; 	// lw
disk[466] <= 32'b000000_00110_00111_10111_00000_000011; 	// div
disk[467] <= 32'b010010_11110_10111_1111111111111111; 	// sw
disk[468] <= 32'b000000_00110_00111_01111_00000_000100; 	// mod
disk[469] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[470] <= 32'b000000_01111_10001_10000_00000_010000; 	// gt
disk[471] <= 32'b010101_10000_00000_0000000111011100; 	// jf
disk[472] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[473] <= 32'b000001_01000_10010_0000000000000001; 	// addi
disk[474] <= 32'b010010_11110_10010_1111111111111111; 	// sw
disk[475] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[476] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[477] <= 32'b010010_11110_10011_1111111111111110; 	// sw
disk[478] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[479] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[480] <= 32'b000000_00101_00110_10100_00000_001110; 	// lt
disk[481] <= 32'b010101_10100_00000_0000000111101010; 	// jf
disk[482] <= 32'b010001_11101_00111_0000000001101011; 	// la
disk[483] <= 32'b000000_00111_00101_10101_00000_000000; 	// add
disk[484] <= 32'b010000_00000_10110_0000000000000001; 	// li
disk[485] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[486] <= 32'b000001_00101_10111_0000000000000001; 	// addi
disk[487] <= 32'b010010_11110_10111_1111111111111110; 	// sw
disk[488] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[489] <= 32'b111100_00000000000000000111011110; 	// j
disk[490] <= 32'b001110_11110_01111_0000000000000000; 	// mov
disk[491] <= 32'b001111_11101_00101_0000000011101011; 	// lw
disk[492] <= 32'b000000_01111_00101_10000_00000_000011; 	// div
disk[493] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[494] <= 32'b001110_11110_10001_0000000000000000; 	// mov
disk[495] <= 32'b000000_10001_00101_10010_00000_000100; 	// mod
disk[496] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[497] <= 32'b000000_10010_10100_10011_00000_010000; 	// gt
disk[498] <= 32'b010101_10011_00000_0000000111110111; 	// jf
disk[499] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[500] <= 32'b000001_00110_10101_0000000000000001; 	// addi
disk[501] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[502] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[503] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[504] <= 32'b000001_00101_10110_0000000000000001; 	// addi
disk[505] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[506] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[507] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[508] <= 32'b010010_11110_10111_1111111111111110; 	// sw
disk[509] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[510] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[511] <= 32'b000000_00101_00110_01111_00000_001110; 	// lt
disk[512] <= 32'b010101_01111_00000_0000001000001001; 	// jf
disk[513] <= 32'b010001_11101_00111_0000000011110100; 	// la
disk[514] <= 32'b000000_00111_00101_10000_00000_000000; 	// add
disk[515] <= 32'b010000_00000_10001_0000000000000001; 	// li
disk[516] <= 32'b010010_10000_10001_0000000000000000; 	// sw
disk[517] <= 32'b000001_00101_10010_0000000000000001; 	// addi
disk[518] <= 32'b010010_11110_10010_1111111111111110; 	// sw
disk[519] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[520] <= 32'b111100_00000000000000000111111101; 	// j
disk[521] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[522] <= 32'b001111_11101_00110_0000000011101011; 	// lw
disk[523] <= 32'b000000_00101_00110_10011_00000_000010; 	// mul
disk[524] <= 32'b010010_11101_10011_0000000011110001; 	// sw
disk[525] <= 32'b001111_11101_00111_0000000011101100; 	// lw
disk[526] <= 32'b000010_00111_10100_0000000000000001; 	// subi
disk[527] <= 32'b010001_11101_01000_0000000011110100; 	// la
disk[528] <= 32'b000000_01000_10100_10101_00000_000000; 	// add
disk[529] <= 32'b010000_00000_10110_0000000000000001; 	// li
disk[530] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[531] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[532] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[533] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[534] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[535] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[536] <= 32'b001111_11101_00110_0000000011101110; 	// lw
disk[537] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[538] <= 32'b010101_10000_00000_0000001000110011; 	// jf
disk[539] <= 32'b010001_11101_00111_0000000101110110; 	// la
disk[540] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[541] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[542] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[543] <= 32'b010001_11101_01000_0000000110000000; 	// la
disk[544] <= 32'b000000_01000_00101_10011_00000_000000; 	// add
disk[545] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[546] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[547] <= 32'b010001_11101_01001_0000000110001010; 	// la
disk[548] <= 32'b000000_01001_00101_10101_00000_000000; 	// add
disk[549] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[550] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[551] <= 32'b010001_11101_01010_0000000110010100; 	// la
disk[552] <= 32'b000000_01010_00101_10111_00000_000000; 	// add
disk[553] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[554] <= 32'b010010_10111_01111_0000000000000000; 	// sw
disk[555] <= 32'b010001_11101_01011_0000000110011110; 	// la
disk[556] <= 32'b000000_01011_00101_10000_00000_000000; 	// add
disk[557] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[558] <= 32'b010010_10000_10001_0000000000000000; 	// sw
disk[559] <= 32'b000001_00101_10010_0000000000000001; 	// addi
disk[560] <= 32'b010010_11110_10010_1111111111111111; 	// sw
disk[561] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[562] <= 32'b111100_00000000000000001000010111; 	// j
disk[563] <= 32'b001111_11101_00101_0000000011101111; 	// lw
disk[564] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[565] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[566] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[567] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[568] <= 32'b001111_11101_00110_0000000011110000; 	// lw
disk[569] <= 32'b000000_00101_00110_10100_00000_001110; 	// lt
disk[570] <= 32'b010101_10100_00000_0000001001011000; 	// jf
disk[571] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[572] <= 32'b010110_00001_10101_0000000000000000; 	// ldk
disk[573] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[574] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[575] <= 32'b001101_00111_10110_0000000000011010; 	// srli
disk[576] <= 32'b001111_11101_01000_0000000110101001; 	// lw
disk[577] <= 32'b000000_10110_01000_10111_00000_001100; 	// eq
disk[578] <= 32'b010101_10111_00000_0000001001010011; 	// jf
disk[579] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[580] <= 32'b000001_01001_01111_0000000000000001; 	// addi
disk[581] <= 32'b010001_11101_01010_0000000101110110; 	// la
disk[582] <= 32'b000000_01010_01001_10000_00000_000000; 	// add
disk[583] <= 32'b010010_10000_01111_0000000000000000; 	// sw
disk[584] <= 32'b000000_01010_01001_10001_00000_000000; 	// add
disk[585] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[586] <= 32'b010001_11101_01011_0000000110001010; 	// la
disk[587] <= 32'b000000_01011_01001_10010_00000_000000; 	// add
disk[588] <= 32'b010010_10010_10001_0000000000000000; 	// sw
disk[589] <= 32'b010001_11101_01100_0000000110000000; 	// la
disk[590] <= 32'b000000_01100_01001_10011_00000_000000; 	// add
disk[591] <= 32'b010010_10011_00101_0000000000000000; 	// sw
disk[592] <= 32'b000001_01001_10100_0000000000000001; 	// addi
disk[593] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[594] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[595] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[596] <= 32'b000001_00101_10101_0000000000000001; 	// addi
disk[597] <= 32'b010010_11110_10101_1111111111111110; 	// sw
disk[598] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[599] <= 32'b111100_00000000000000001000110111; 	// j
disk[600] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[601] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[602] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[603] <= 32'b111110_00000000000000000101001011; 	// jal
disk[604] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[605] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[606] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[607] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[608] <= 32'b111110_00000000000000000110000101; 	// jal
disk[609] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[610] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[611] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[612] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[613] <= 32'b111110_00000000000000000110010001; 	// jal
disk[614] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[615] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[616] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[617] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[618] <= 32'b111110_00000000000000000110101011; 	// jal
disk[619] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[620] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[621] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[622] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[623] <= 32'b111110_00000000000000000110110101; 	// jal
disk[624] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[625] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[626] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[627] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[628] <= 32'b111110_00000000000000001000010100; 	// jal
disk[629] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[630] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[631] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[632] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[633] <= 32'b111110_00000000000000000101000101; 	// jal
disk[634] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[635] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[636] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[637] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[638] <= 32'b000001_11110_11110_0000000000000110; 	// addi
disk[639] <= 32'b010010_11110_00001_1111111111111101; 	// sw
disk[640] <= 32'b001111_11110_00101_1111111111111101; 	// lw
disk[641] <= 32'b001111_11101_00110_0000000011101011; 	// lw
disk[642] <= 32'b000000_00101_00110_01111_00000_000011; 	// div
disk[643] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[644] <= 32'b000000_00101_00110_10000_00000_000100; 	// mod
disk[645] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[646] <= 32'b000000_10000_10010_10001_00000_010000; 	// gt
disk[647] <= 32'b010101_10001_00000_0000001010001100; 	// jf
disk[648] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[649] <= 32'b000001_00111_10011_0000000000000001; 	// addi
disk[650] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[651] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[652] <= 32'b010001_11101_00101_0000000001001010; 	// la
disk[653] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[654] <= 32'b000000_00101_00110_10100_00000_000000; 	// add
disk[655] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[656] <= 32'b010010_10100_00111_0000000000000000; 	// sw
disk[657] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[658] <= 32'b010010_11110_10101_1111111111111110; 	// sw
disk[659] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[660] <= 32'b001111_11101_00110_0000000011101100; 	// lw
disk[661] <= 32'b000000_00101_00110_10110_00000_001110; 	// lt
disk[662] <= 32'b010101_10110_00000_0000001010110110; 	// jf
disk[663] <= 32'b010001_11101_00111_0000000001101011; 	// la
disk[664] <= 32'b000000_00111_00101_10111_00000_000000; 	// add
disk[665] <= 32'b001111_10111_10111_0000000000000000; 	// lw
disk[666] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[667] <= 32'b000000_10111_10000_01111_00000_001100; 	// eq
disk[668] <= 32'b010101_01111_00000_0000001010110001; 	// jf
disk[669] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[670] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[671] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[672] <= 32'b000000_00101_10010_10001_00000_010000; 	// gt
disk[673] <= 32'b010101_10001_00000_0000001010101110; 	// jf
disk[674] <= 32'b010001_11101_00110_0000000001101011; 	// la
disk[675] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[676] <= 32'b000000_00110_00111_10011_00000_000000; 	// add
disk[677] <= 32'b010000_00000_10100_0000000000000001; 	// li
disk[678] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[679] <= 32'b000010_00101_10101_0000000000000001; 	// subi
disk[680] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[681] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[682] <= 32'b000001_00111_10110_0000000000000001; 	// addi
disk[683] <= 32'b010010_11110_10110_1111111111111110; 	// sw
disk[684] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[685] <= 32'b111100_00000000000000001010011110; 	// j
disk[686] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[687] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[688] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[689] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[690] <= 32'b000001_00101_10111_0000000000000001; 	// addi
disk[691] <= 32'b010010_11110_10111_1111111111111110; 	// sw
disk[692] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[693] <= 32'b111100_00000000000000001010010011; 	// j
disk[694] <= 32'b001111_11101_00101_0000000011101101; 	// lw
disk[695] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[696] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[697] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[698] <= 32'b010001_11101_00101_0000000000011000; 	// la
disk[699] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[700] <= 32'b000000_00101_00110_01111_00000_000000; 	// add
disk[701] <= 32'b001111_01111_01111_0000000000000000; 	// lw
disk[702] <= 32'b001111_11101_00111_0000000011101011; 	// lw
disk[703] <= 32'b000000_01111_00111_10000_00000_000011; 	// div
disk[704] <= 32'b000001_10000_10001_0000000000000001; 	// addi
disk[705] <= 32'b010010_11110_10001_1111111111111111; 	// sw
disk[706] <= 32'b000000_00101_00110_10010_00000_000000; 	// add
disk[707] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[708] <= 32'b000000_10010_00111_10011_00000_000100; 	// mod
disk[709] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[710] <= 32'b000000_10011_10101_10100_00000_010000; 	// gt
disk[711] <= 32'b010101_10100_00000_0000001011001100; 	// jf
disk[712] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[713] <= 32'b000001_01000_10110_0000000000000001; 	// addi
disk[714] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[715] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[716] <= 32'b001111_11101_00101_0000000011101100; 	// lw
disk[717] <= 32'b000010_00101_10111_0000000000000001; 	// subi
disk[718] <= 32'b010010_11110_10111_1111111111111110; 	// sw
disk[719] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[720] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[721] <= 32'b000000_00101_10000_01111_00000_010000; 	// gt
disk[722] <= 32'b010101_01111_00000_0000001011110010; 	// jf
disk[723] <= 32'b010001_11101_00110_0000000011110100; 	// la
disk[724] <= 32'b000000_00110_00101_10001_00000_000000; 	// add
disk[725] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[726] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[727] <= 32'b000000_10001_10011_10010_00000_001100; 	// eq
disk[728] <= 32'b010101_10010_00000_0000001011101101; 	// jf
disk[729] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[730] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[731] <= 32'b000000_00101_10101_10100_00000_010000; 	// gt
disk[732] <= 32'b010101_10100_00000_0000001011101010; 	// jf
disk[733] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[734] <= 32'b010010_11110_00110_0000000000000000; 	// sw
disk[735] <= 32'b010001_11101_00111_0000000011110100; 	// la
disk[736] <= 32'b000000_00111_00110_10110_00000_000000; 	// add
disk[737] <= 32'b010000_00000_10111_0000000000000001; 	// li
disk[738] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[739] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[740] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[741] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[742] <= 32'b000010_00110_10000_0000000000000001; 	// subi
disk[743] <= 32'b010010_11110_10000_1111111111111110; 	// sw
disk[744] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[745] <= 32'b111100_00000000000000001011011001; 	// j
disk[746] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[747] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[748] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[749] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[750] <= 32'b000010_00101_10001_0000000000000001; 	// subi
disk[751] <= 32'b010010_11110_10001_1111111111111110; 	// sw
disk[752] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[753] <= 32'b111100_00000000000000001011001111; 	// j
disk[754] <= 32'b001111_11101_00101_0000000011101101; 	// lw
disk[755] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[756] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[757] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[758] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[759] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[760] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[761] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[762] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[763] <= 32'b001111_11101_00110_0000000011101110; 	// lw
disk[764] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[765] <= 32'b010101_10001_00000_0000001100010011; 	// jf
disk[766] <= 32'b010001_11101_00111_0000000110010100; 	// la
disk[767] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
disk[768] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[769] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[770] <= 32'b000000_10010_10100_10011_00000_001101; 	// ne
disk[771] <= 32'b010101_10011_00000_0000001100001110; 	// jf
disk[772] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[773] <= 32'b010010_11110_11111_1111111111111110; 	// sw
disk[774] <= 32'b111110_00000000000000000000011001; 	// jal
disk[775] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[776] <= 32'b001111_11110_11111_1111111111111110; 	// lw
disk[777] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[778] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[779] <= 32'b000000_00110_00101_10101_00000_000000; 	// add
disk[780] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[781] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[782] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[783] <= 32'b000001_00101_10110_0000000000000001; 	// addi
disk[784] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[785] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[786] <= 32'b111100_00000000000000001011111010; 	// j
disk[787] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[788] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[789] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[790] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[791] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[792] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[793] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[794] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[795] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[796] <= 32'b001111_11101_00110_0000000011101110; 	// lw
disk[797] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[798] <= 32'b010101_10001_00000_0000001100110100; 	// jf
disk[799] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[800] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
disk[801] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[802] <= 32'b001111_11101_01000_0000000000000010; 	// lw
disk[803] <= 32'b000000_10010_01000_10011_00000_001100; 	// eq
disk[804] <= 32'b010101_10011_00000_0000001100101111; 	// jf
disk[805] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[806] <= 32'b010010_11110_11111_1111111111111110; 	// sw
disk[807] <= 32'b111110_00000000000000000000011001; 	// jal
disk[808] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[809] <= 32'b001111_11110_11111_1111111111111110; 	// lw
disk[810] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[811] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[812] <= 32'b000000_00110_00101_10100_00000_000000; 	// add
disk[813] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[814] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[815] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[816] <= 32'b000001_00101_10101_0000000000000001; 	// addi
disk[817] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[818] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[819] <= 32'b111100_00000000000000001100011011; 	// j
disk[820] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[821] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[822] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[823] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[824] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[825] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[826] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[827] <= 32'b001111_11101_00110_0000000011101110; 	// lw
disk[828] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[829] <= 32'b010101_10000_00000_0000001101001011; 	// jf
disk[830] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[831] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[832] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[833] <= 32'b001111_11101_01000_0000000000000010; 	// lw
disk[834] <= 32'b000000_10001_01000_10010_00000_001100; 	// eq
disk[835] <= 32'b010101_10010_00000_0000001101000110; 	// jf
disk[836] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[837] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[838] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[839] <= 32'b000001_00101_10011_0000000000000001; 	// addi
disk[840] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[841] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[842] <= 32'b111100_00000000000000001100111010; 	// j
disk[843] <= 32'b001111_11101_00101_0000000000000011; 	// lw
disk[844] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[845] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[846] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[847] <= 32'b010010_11110_00001_1111111111111110; 	// sw
disk[848] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[849] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[850] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[851] <= 32'b001111_11101_00110_0000000011101110; 	// lw
disk[852] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[853] <= 32'b010101_10000_00000_0000001101100110; 	// jf
disk[854] <= 32'b010001_11101_00111_0000000001100000; 	// la
disk[855] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[856] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[857] <= 32'b001111_11110_01000_1111111111111110; 	// lw
disk[858] <= 32'b000000_10001_01000_10010_00000_001100; 	// eq
disk[859] <= 32'b010101_10010_00000_0000001101100001; 	// jf
disk[860] <= 32'b000000_00111_00101_10011_00000_000000; 	// add
disk[861] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[862] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[863] <= 32'b000001_00101_10101_0000000000000001; 	// addi
disk[864] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[865] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[866] <= 32'b000001_00101_10110_0000000000000001; 	// addi
disk[867] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[868] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[869] <= 32'b111100_00000000000000001101010010; 	// j
disk[870] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[871] <= 32'b001111_11101_00110_0000000011101110; 	// lw
disk[872] <= 32'b000000_00101_00110_10111_00000_001110; 	// lt
disk[873] <= 32'b010101_10111_00000_0000001101110100; 	// jf
disk[874] <= 32'b010001_11101_00111_0000000001100000; 	// la
disk[875] <= 32'b000000_00111_00101_01111_00000_000000; 	// add
disk[876] <= 32'b001111_01111_01111_0000000000000000; 	// lw
disk[877] <= 32'b000010_00101_10000_0000000000000001; 	// subi
disk[878] <= 32'b000000_00111_10000_10001_00000_000000; 	// add
disk[879] <= 32'b010010_10001_01111_0000000000000000; 	// sw
disk[880] <= 32'b000001_00101_10010_0000000000000001; 	// addi
disk[881] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[882] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[883] <= 32'b111100_00000000000000001101100110; 	// j
disk[884] <= 32'b001111_11101_00101_0000000011101110; 	// lw
disk[885] <= 32'b000010_00101_10011_0000000000000001; 	// subi
disk[886] <= 32'b010001_11101_00110_0000000001100000; 	// la
disk[887] <= 32'b000000_00110_10011_10100_00000_000000; 	// add
disk[888] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[889] <= 32'b010010_10100_10101_0000000000000000; 	// sw
disk[890] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[891] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[892] <= 32'b010000_00000_01111_0000000000000001; 	// li
disk[893] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[894] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[895] <= 32'b001111_11101_00110_0000000011101110; 	// lw
disk[896] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[897] <= 32'b010101_10000_00000_0000001110001100; 	// jf
disk[898] <= 32'b010001_11101_00111_0000000001100000; 	// la
disk[899] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[900] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[901] <= 32'b000010_00101_10010_0000000000000001; 	// subi
disk[902] <= 32'b000000_00111_10010_10011_00000_000000; 	// add
disk[903] <= 32'b010010_10011_10001_0000000000000000; 	// sw
disk[904] <= 32'b000001_00101_10100_0000000000000001; 	// addi
disk[905] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[906] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[907] <= 32'b111100_00000000000000001101111110; 	// j
disk[908] <= 32'b001111_11101_00101_0000000011101110; 	// lw
disk[909] <= 32'b000010_00101_10101_0000000000000001; 	// subi
disk[910] <= 32'b010001_11101_00110_0000000001100000; 	// la
disk[911] <= 32'b000000_00110_10101_10110_00000_000000; 	// add
disk[912] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[913] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[914] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[915] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[916] <= 32'b010001_11101_00101_0000000001100000; 	// la
disk[917] <= 32'b001111_00101_01111_0000000000000000; 	// lw
disk[918] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[919] <= 32'b000000_01111_10001_10000_00000_001101; 	// ne
disk[920] <= 32'b010101_10000_00000_0000001110100011; 	// jf
disk[921] <= 32'b001111_00101_10010_0000000000000000; 	// lw
disk[922] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[923] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[924] <= 32'b111110_00000000000000001101111011; 	// jal
disk[925] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[926] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[927] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[928] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[929] <= 32'b001110_00110_11000_0000000000000000; 	// mov
disk[930] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[931] <= 32'b001111_11101_00101_0000000000000011; 	// lw
disk[932] <= 32'b001110_00101_11000_0000000000000000; 	// mov
disk[933] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[934] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[935] <= 32'b010010_11110_00001_1111111111111111; 	// sw
disk[936] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[937] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[938] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[939] <= 32'b001111_11101_00110_0000000011101110; 	// lw
disk[940] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[941] <= 32'b010101_10000_00000_0000001110111101; 	// jf
disk[942] <= 32'b010001_11101_00111_0000000001100000; 	// la
disk[943] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[944] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[945] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[946] <= 32'b000000_10001_10011_10010_00000_001100; 	// eq
disk[947] <= 32'b010101_10010_00000_0000001110111000; 	// jf
disk[948] <= 32'b000000_00111_00101_10100_00000_000000; 	// add
disk[949] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[950] <= 32'b010010_10100_01000_0000000000000000; 	// sw
disk[951] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[952] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[953] <= 32'b000001_00101_10101_0000000000000001; 	// addi
disk[954] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[955] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[956] <= 32'b111100_00000000000000001110101010; 	// j
disk[957] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[958] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[959] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[960] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[961] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[962] <= 32'b001111_11101_00110_0000000011101110; 	// lw
disk[963] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[964] <= 32'b010101_10000_00000_0000001111100000; 	// jf
disk[965] <= 32'b010001_11101_00111_0000000110010100; 	// la
disk[966] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[967] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[968] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[969] <= 32'b000000_10001_10011_10010_00000_001101; 	// ne
disk[970] <= 32'b010101_10010_00000_0000001111011011; 	// jf
disk[971] <= 32'b010001_11101_01000_0000000000000100; 	// la
disk[972] <= 32'b000000_01000_00101_10100_00000_000000; 	// add
disk[973] <= 32'b001111_10100_10100_0000000000000000; 	// lw
disk[974] <= 32'b001111_11101_01001_0000000000000010; 	// lw
disk[975] <= 32'b000000_10100_01001_10101_00000_001101; 	// ne
disk[976] <= 32'b010101_10101_00000_0000001111011011; 	// jf
disk[977] <= 32'b000000_01000_00101_10110_00000_000000; 	// add
disk[978] <= 32'b001111_11101_01010_0000000000000001; 	// lw
disk[979] <= 32'b010010_10110_01010_0000000000000000; 	// sw
disk[980] <= 32'b000001_00101_10111_0000000000000001; 	// addi
disk[981] <= 32'b001110_10111_00001_0000000000000000; 	// mov
disk[982] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[983] <= 32'b111110_00000000000000001110100110; 	// jal
disk[984] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[985] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[986] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[987] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[988] <= 32'b000001_00101_01111_0000000000000001; 	// addi
disk[989] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[990] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[991] <= 32'b111100_00000000000000001111000001; 	// j
disk[992] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[993] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[994] <= 32'b010010_11110_00001_1111111111111110; 	// sw
disk[995] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[996] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[997] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[998] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[999] <= 32'b010110_00001_01111_0000000000000000; 	// ldk
disk[1000] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[1001] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[1002] <= 32'b001101_00101_10000_0000000000011010; 	// srli
disk[1003] <= 32'b001111_11101_00110_0000000110101000; 	// lw
disk[1004] <= 32'b000000_10000_00110_10001_00000_001101; 	// ne
disk[1005] <= 32'b010101_10001_00000_0000001111110111; 	// jf
disk[1006] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[1007] <= 32'b000001_00111_10010_0000000000000001; 	// addi
disk[1008] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[1009] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[1010] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1011] <= 32'b010110_00001_10011_0000000000000000; 	// ldk
disk[1012] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[1013] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[1014] <= 32'b111100_00000000000000001111101001; 	// j
disk[1015] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1016] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[1017] <= 32'b000000_00101_00110_10100_00000_000001; 	// sub
disk[1018] <= 32'b001110_10100_11000_0000000000000000; 	// mov
disk[1019] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[1020] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[1021] <= 32'b010010_11110_00001_1111111111111111; 	// sw
disk[1022] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[1023] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[1024] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1025] <= 32'b001111_11101_00110_0000000011101110; 	// lw
disk[1026] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[1027] <= 32'b010101_10000_00000_0000010000010101; 	// jf
disk[1028] <= 32'b010001_11101_00111_0000000110001010; 	// la
disk[1029] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[1030] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[1031] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[1032] <= 32'b000000_10001_01000_10010_00000_001100; 	// eq
disk[1033] <= 32'b010101_10010_00000_0000010000010000; 	// jf
disk[1034] <= 32'b010001_11101_01001_0000000101110110; 	// la
disk[1035] <= 32'b000000_01001_00101_10011_00000_000000; 	// add
disk[1036] <= 32'b001111_10011_10011_0000000000000000; 	// lw
disk[1037] <= 32'b000010_10011_10100_0000000000000001; 	// subi
disk[1038] <= 32'b001110_10100_11000_0000000000000000; 	// mov
disk[1039] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[1040] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1041] <= 32'b000001_00101_10101_0000000000000001; 	// addi
disk[1042] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[1043] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1044] <= 32'b111100_00000000000000010000000000; 	// j
disk[1045] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[1046] <= 32'b000001_11110_11110_0000000000001010; 	// addi
disk[1047] <= 32'b010010_11110_00001_1111111111111001; 	// sw
disk[1048] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1049] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1050] <= 32'b010010_11110_11111_1111111111111000; 	// sw
disk[1051] <= 32'b111110_00000000000000001111111100; 	// jal
disk[1052] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1053] <= 32'b001111_11110_11111_1111111111111000; 	// lw
disk[1054] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1055] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1056] <= 32'b001111_11110_00110_1111111111111001; 	// lw
disk[1057] <= 32'b010010_11101_00110_0000000001011111; 	// sw
disk[1058] <= 32'b010001_11101_00111_0000000110000000; 	// la
disk[1059] <= 32'b000000_00111_00110_01111_00000_000000; 	// add
disk[1060] <= 32'b001111_01111_01111_0000000000000000; 	// lw
disk[1061] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[1062] <= 32'b010001_11101_01000_0000000101110110; 	// la
disk[1063] <= 32'b000000_01000_00110_10000_00000_000000; 	// add
disk[1064] <= 32'b001111_10000_10000_0000000000000000; 	// lw
disk[1065] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[1066] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[1067] <= 32'b010010_11110_01001_1111111111111010; 	// sw
disk[1068] <= 32'b001110_01001_00001_0000000000000000; 	// mov
disk[1069] <= 32'b010010_11110_11111_1111111111111000; 	// sw
disk[1070] <= 32'b111110_00000000000000001111100001; 	// jal
disk[1071] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[1072] <= 32'b001111_11110_11111_1111111111111000; 	// lw
disk[1073] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1074] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[1075] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[1076] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1077] <= 32'b010010_11110_11111_1111111111111000; 	// sw
disk[1078] <= 32'b111110_00000000000000001001111110; 	// jal
disk[1079] <= 32'b000010_11110_11110_0000000000000110; 	// subi
disk[1080] <= 32'b001111_11110_11111_1111111111111000; 	// lw
disk[1081] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1082] <= 32'b010010_11110_00101_1111111111111101; 	// sw
disk[1083] <= 32'b010001_11101_00110_0000000000110110; 	// la
disk[1084] <= 32'b001111_11101_00111_0000000001011111; 	// lw
disk[1085] <= 32'b000000_00110_00111_10001_00000_000000; 	// add
disk[1086] <= 32'b001111_11110_01000_1111111111111101; 	// lw
disk[1087] <= 32'b010010_10001_01000_0000000000000000; 	// sw
disk[1088] <= 32'b001111_11101_01001_0000000011101011; 	// lw
disk[1089] <= 32'b000000_01001_01000_10010_00000_000010; 	// mul
disk[1090] <= 32'b010010_11110_10010_1111111111111011; 	// sw
disk[1091] <= 32'b001111_11110_01010_1111111111111010; 	// lw
disk[1092] <= 32'b001110_01010_00001_0000000000000000; 	// mov
disk[1093] <= 32'b010110_00001_10011_0000000000000000; 	// ldk
disk[1094] <= 32'b010010_11110_10011_1111111111111100; 	// sw
disk[1095] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[1096] <= 32'b001101_00101_10100_0000000000011010; 	// srli
disk[1097] <= 32'b001111_11101_00110_0000000110101000; 	// lw
disk[1098] <= 32'b000000_10100_00110_10101_00000_001101; 	// ne
disk[1099] <= 32'b010101_10101_00000_0000010001011100; 	// jf
disk[1100] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1101] <= 32'b001111_11110_00111_1111111111111011; 	// lw
disk[1102] <= 32'b001110_00111_00010_0000000000000000; 	// mov
disk[1103] <= 32'b011001_00010_00001_0000000000000000; 	// sim
disk[1104] <= 32'b001111_11110_01000_1111111111111010; 	// lw
disk[1105] <= 32'b000001_01000_10110_0000000000000001; 	// addi
disk[1106] <= 32'b010010_11110_10110_1111111111111010; 	// sw
disk[1107] <= 32'b001111_11110_01000_1111111111111010; 	// lw
disk[1108] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[1109] <= 32'b010110_00001_10111_0000000000000000; 	// ldk
disk[1110] <= 32'b010010_11110_10111_1111111111111100; 	// sw
disk[1111] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[1112] <= 32'b000001_00111_01111_0000000000000001; 	// addi
disk[1113] <= 32'b010010_11110_01111_1111111111111011; 	// sw
disk[1114] <= 32'b001111_11110_00111_1111111111111011; 	// lw
disk[1115] <= 32'b111100_00000000000000010001000111; 	// j
disk[1116] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[1117] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1118] <= 32'b001111_11110_00110_1111111111111011; 	// lw
disk[1119] <= 32'b001110_00110_00010_0000000000000000; 	// mov
disk[1120] <= 32'b011001_00010_00001_0000000000000000; 	// sim
disk[1121] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[1122] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1123] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
disk[1124] <= 32'b001111_11101_01000_0000000011101011; 	// lw
disk[1125] <= 32'b001111_11110_01001_1111111111111101; 	// lw
disk[1126] <= 32'b000000_01000_01001_10000_00000_000010; 	// mul
disk[1127] <= 32'b001110_10000_00001_0000000000000000; 	// mov
disk[1128] <= 32'b011010_00000_00001_0000000000000000; 	// mmuLowerIM
disk[1129] <= 32'b010001_11101_01010_0000000110010100; 	// la
disk[1130] <= 32'b001111_11110_01011_1111111111111001; 	// lw
disk[1131] <= 32'b000000_01010_01011_10001_00000_000000; 	// add
disk[1132] <= 32'b010010_10001_00111_0000000000000000; 	// sw
disk[1133] <= 32'b010001_11101_01100_0000000110011110; 	// la
disk[1134] <= 32'b000000_01100_01011_10010_00000_000000; 	// add
disk[1135] <= 32'b001111_11110_01101_1111111111111111; 	// lw
disk[1136] <= 32'b010010_10010_01101_0000000000000000; 	// sw
disk[1137] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[1138] <= 32'b010010_11101_10011_0000000001011111; 	// sw
disk[1139] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[1140] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[1141] <= 32'b010010_11110_00001_0000000000000000; 	// sw
disk[1142] <= 32'b010001_11101_00101_0000000110010100; 	// la
disk[1143] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[1144] <= 32'b000000_00101_00110_01111_00000_000000; 	// add
disk[1145] <= 32'b001111_01111_01111_0000000000000000; 	// lw
disk[1146] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[1147] <= 32'b000000_01111_10001_10000_00000_001101; 	// ne
disk[1148] <= 32'b010101_10000_00000_0000010010101000; 	// jf
disk[1149] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[1150] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1151] <= 32'b100100_00000_00001_0000000000000000; 	// lcdCurr
disk[1152] <= 32'b001111_11101_01000_0000000110110101; 	// lw
disk[1153] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[1154] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[1155] <= 32'b001111_11101_01001_0000000011110001; 	// lw
disk[1156] <= 32'b000001_01001_10010_0000000000000001; 	// addi
disk[1157] <= 32'b010010_11101_10010_0000000011110010; 	// sw
disk[1158] <= 32'b010001_11101_01010_0000000000000100; 	// la
disk[1159] <= 32'b000000_01010_00110_10011_00000_000000; 	// add
disk[1160] <= 32'b001111_11101_01011_0000000000000000; 	// lw
disk[1161] <= 32'b010010_10011_01011_0000000000000000; 	// sw
disk[1162] <= 32'b010001_11101_01100_0000000000001110; 	// la
disk[1163] <= 32'b000000_01100_00110_10100_00000_000000; 	// add
disk[1164] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[1165] <= 32'b010010_10100_10101_0000000000000000; 	// sw
disk[1166] <= 32'b001111_11101_01101_0000000011110010; 	// lw
disk[1167] <= 32'b001110_01101_00001_0000000000000000; 	// mov
disk[1168] <= 32'b001110_00001_11100_0000000000000000; 	// mov
disk[1169] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1170] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
disk[1171] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[1172] <= 32'b001110_11110_00011_0000000000000000; 	// mov
disk[1173] <= 32'b001110_11101_00100_0000000000000000; 	// mov
disk[1174] <= 32'b001110_11100_11110_0000000000000000; 	// mov
disk[1175] <= 32'b001110_11011_11101_0000000000000000; 	// mov
disk[1176] <= 32'b001110_00011_11100_0000000000000000; 	// mov
disk[1177] <= 32'b001110_00100_11011_0000000000000000; 	// mov
disk[1178] <= 32'b100000_00000000000000000000000000; 	// exec
disk[1179] <= 32'b001110_11100_11110_0000000000000000; 	// mov
disk[1180] <= 32'b001110_11011_11101_0000000000000000; 	// mov
disk[1181] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[1182] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1183] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1184] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[1185] <= 32'b111110_00000000000000000010000110; 	// jal
disk[1186] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[1187] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[1188] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1189] <= 32'b001111_11101_00110_0000000110101011; 	// lw
disk[1190] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1191] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[1192] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[1193] <= 32'b000001_11110_11110_0000000000001000; 	// addi
disk[1194] <= 32'b010010_11110_00001_1111111111111011; 	// sw
disk[1195] <= 32'b001111_11110_00101_1111111111111011; 	// lw
disk[1196] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1197] <= 32'b100100_00000_00001_0000000000000000; 	// lcdCurr
disk[1198] <= 32'b001111_11101_00110_0000000110110101; 	// lw
disk[1199] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1200] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[1201] <= 32'b001111_11101_00111_0000000011110001; 	// lw
disk[1202] <= 32'b000001_00111_01111_0000000000000001; 	// addi
disk[1203] <= 32'b010010_11101_01111_0000000011110010; 	// sw
disk[1204] <= 32'b010001_11101_01000_0000000000000100; 	// la
disk[1205] <= 32'b001111_11101_01001_0000000001011111; 	// lw
disk[1206] <= 32'b000000_01000_01001_10000_00000_000000; 	// add
disk[1207] <= 32'b001111_11101_01010_0000000000000000; 	// lw
disk[1208] <= 32'b010010_10000_01010_0000000000000000; 	// sw
disk[1209] <= 32'b010001_11101_01011_0000000001000000; 	// la
disk[1210] <= 32'b000000_01011_01001_10001_00000_000000; 	// add
disk[1211] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[1212] <= 32'b010010_11110_10001_1111111111111101; 	// sw
disk[1213] <= 32'b001111_11101_01100_0000000011110010; 	// lw
disk[1214] <= 32'b010010_11110_01100_1111111111111110; 	// sw
disk[1215] <= 32'b001111_11110_01101_1111111111111101; 	// lw
disk[1216] <= 32'b001111_11101_01110_0000000011101011; 	// lw
disk[1217] <= 32'b000000_01101_01110_10010_00000_000010; 	// mul
disk[1218] <= 32'b010010_11110_10010_1111111111111111; 	// sw
disk[1219] <= 32'b010001_11101_00101_0000000000011000; 	// la
disk[1220] <= 32'b000000_00101_01001_10011_00000_000000; 	// add
disk[1221] <= 32'b001111_10011_10011_0000000000000000; 	// lw
disk[1222] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[1223] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1224] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[1225] <= 32'b000000_00101_10101_10100_00000_010000; 	// gt
disk[1226] <= 32'b010101_10100_00000_0000010011011110; 	// jf
disk[1227] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[1228] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1229] <= 32'b001111_00001_10110_0000000000000000; 	// lw
disk[1230] <= 32'b010010_11110_10110_1111111111111100; 	// sw
disk[1231] <= 32'b001111_11110_00111_1111111111111100; 	// lw
disk[1232] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1233] <= 32'b001111_11110_01000_1111111111111110; 	// lw
disk[1234] <= 32'b001110_01000_00010_0000000000000000; 	// mov
disk[1235] <= 32'b010010_00010_00001_0000000000000000; 	// sw
disk[1236] <= 32'b000001_01000_10111_0000000000000001; 	// addi
disk[1237] <= 32'b010010_11110_10111_1111111111111110; 	// sw
disk[1238] <= 32'b001111_11110_01000_1111111111111110; 	// lw
disk[1239] <= 32'b000001_00110_01111_0000000000000001; 	// addi
disk[1240] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[1241] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[1242] <= 32'b000010_00101_10000_0000000000000001; 	// subi
disk[1243] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[1244] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1245] <= 32'b111100_00000000000000010011000111; 	// j
disk[1246] <= 32'b010001_11101_00101_0000000000011000; 	// la
disk[1247] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[1248] <= 32'b000000_00101_00110_10001_00000_000000; 	// add
disk[1249] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[1250] <= 32'b001111_11101_00111_0000000011110001; 	// lw
disk[1251] <= 32'b000000_00111_10001_10010_00000_000000; 	// add
disk[1252] <= 32'b001110_10010_00001_0000000000000000; 	// mov
disk[1253] <= 32'b001110_00001_11100_0000000000000000; 	// mov
disk[1254] <= 32'b000001_00110_10011_0000000000000001; 	// addi
disk[1255] <= 32'b001110_10011_00001_0000000000000000; 	// mov
disk[1256] <= 32'b010001_11101_01000_0000000000001110; 	// la
disk[1257] <= 32'b000000_01000_00110_10100_00000_000000; 	// add
disk[1258] <= 32'b001111_10100_10100_0000000000000000; 	// lw
disk[1259] <= 32'b001110_10100_00010_0000000000000000; 	// mov
disk[1260] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
disk[1261] <= 32'b010010_11110_11111_1111111111111010; 	// sw
disk[1262] <= 32'b001110_11110_00011_0000000000000000; 	// mov
disk[1263] <= 32'b001110_11101_00100_0000000000000000; 	// mov
disk[1264] <= 32'b001110_11100_11110_0000000000000000; 	// mov
disk[1265] <= 32'b001110_11011_11101_0000000000000000; 	// mov
disk[1266] <= 32'b001110_00011_11100_0000000000000000; 	// mov
disk[1267] <= 32'b001110_00100_11011_0000000000000000; 	// mov
disk[1268] <= 32'b001110_00010_11010_0000000000000000; 	// mov
disk[1269] <= 32'b001111_00000_00000_0000111111100000; 	// lw
disk[1270] <= 32'b001111_00000_00001_0000111111100001; 	// lw
disk[1271] <= 32'b001111_00000_00010_0000111111100010; 	// lw
disk[1272] <= 32'b001111_00000_00011_0000111111100011; 	// lw
disk[1273] <= 32'b001111_00000_00100_0000111111100100; 	// lw
disk[1274] <= 32'b001111_00000_00101_0000111111100101; 	// lw
disk[1275] <= 32'b001111_00000_00110_0000111111100110; 	// lw
disk[1276] <= 32'b001111_00000_00111_0000111111100111; 	// lw
disk[1277] <= 32'b001111_00000_01000_0000111111101000; 	// lw
disk[1278] <= 32'b001111_00000_01001_0000111111101001; 	// lw
disk[1279] <= 32'b001111_00000_01010_0000111111101010; 	// lw
disk[1280] <= 32'b001111_00000_01011_0000111111101011; 	// lw
disk[1281] <= 32'b001111_00000_01100_0000111111101100; 	// lw
disk[1282] <= 32'b001111_00000_01101_0000111111101101; 	// lw
disk[1283] <= 32'b001111_00000_01110_0000111111101110; 	// lw
disk[1284] <= 32'b001111_00000_01111_0000111111101111; 	// lw
disk[1285] <= 32'b001111_00000_10000_0000111111110000; 	// lw
disk[1286] <= 32'b001111_00000_10001_0000111111110001; 	// lw
disk[1287] <= 32'b001111_00000_10010_0000111111110010; 	// lw
disk[1288] <= 32'b001111_00000_10011_0000111111110011; 	// lw
disk[1289] <= 32'b001111_00000_10100_0000111111110100; 	// lw
disk[1290] <= 32'b001111_00000_10101_0000111111110101; 	// lw
disk[1291] <= 32'b001111_00000_10110_0000111111110110; 	// lw
disk[1292] <= 32'b001111_00000_10111_0000111111110111; 	// lw
disk[1293] <= 32'b001111_00000_11000_0000111111111000; 	// lw
disk[1294] <= 32'b001111_00000_11111_0000111111111001; 	// lw
disk[1295] <= 32'b100001_11010_00000_0000000000000000; 	// execAgain
disk[1296] <= 32'b001110_11100_11110_0000000000000000; 	// mov
disk[1297] <= 32'b001110_11011_11101_0000000000000000; 	// mov
disk[1298] <= 32'b001111_11110_11111_1111111111111010; 	// lw
disk[1299] <= 32'b001111_11110_00101_1111111111111011; 	// lw
disk[1300] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1301] <= 32'b010010_11110_11111_1111111111111010; 	// sw
disk[1302] <= 32'b111110_00000000000000000010000110; 	// jal
disk[1303] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[1304] <= 32'b001111_11110_11111_1111111111111010; 	// lw
disk[1305] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1306] <= 32'b001111_11101_00110_0000000110101011; 	// lw
disk[1307] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1308] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[1309] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[1310] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[1311] <= 32'b010010_11110_00001_0000000000000000; 	// sw
disk[1312] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1313] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[1314] <= 32'b010010_11101_01111_0000000001011111; 	// sw
disk[1315] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[1316] <= 32'b010010_11101_00110_0000000001011110; 	// sw
disk[1317] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[1318] <= 32'b111110_00000000000000000000111110; 	// jal
disk[1319] <= 32'b000010_11110_11110_0000000000000110; 	// subi
disk[1320] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[1321] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1322] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[1323] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1324] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[1325] <= 32'b111110_00000000000000010010101001; 	// jal
disk[1326] <= 32'b000010_11110_11110_0000000000001000; 	// subi
disk[1327] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[1328] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1329] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[1330] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[1331] <= 32'b010010_11110_00001_0000000000000000; 	// sw
disk[1332] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1333] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[1334] <= 32'b010010_11101_01111_0000000001011111; 	// sw
disk[1335] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[1336] <= 32'b010010_11101_00110_0000000001011110; 	// sw
disk[1337] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1338] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[1339] <= 32'b111110_00000000000000010001110100; 	// jal
disk[1340] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1341] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[1342] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1343] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[1344] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[1345] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[1346] <= 32'b111110_00000000000000001110111110; 	// jal
disk[1347] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1348] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[1349] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1350] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[1351] <= 32'b111110_00000000000000001110010011; 	// jal
disk[1352] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1353] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[1354] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1355] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[1356] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1357] <= 32'b001111_11101_00110_0000000000000011; 	// lw
disk[1358] <= 32'b000000_00101_00110_01111_00000_001101; 	// ne
disk[1359] <= 32'b010101_01111_00000_0000010101110011; 	// jf
disk[1360] <= 32'b000010_00101_10000_0000000000000001; 	// subi
disk[1361] <= 32'b010010_11101_10000_0000000001011111; 	// sw
disk[1362] <= 32'b010001_11101_00111_0000000000001110; 	// la
disk[1363] <= 32'b001111_11101_01000_0000000001011111; 	// lw
disk[1364] <= 32'b000000_00111_01000_10001_00000_000000; 	// add
disk[1365] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[1366] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[1367] <= 32'b000000_10001_10011_10010_00000_001100; 	// eq
disk[1368] <= 32'b010101_10010_00000_0000010101100000; 	// jf
disk[1369] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1370] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[1371] <= 32'b111110_00000000000000010001110100; 	// jal
disk[1372] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1373] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[1374] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1375] <= 32'b111100_00000000000000010101101100; 	// j
disk[1376] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[1377] <= 32'b111110_00000000000000000000111110; 	// jal
disk[1378] <= 32'b000010_11110_11110_0000000000000110; 	// subi
disk[1379] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[1380] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1381] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[1382] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1383] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[1384] <= 32'b111110_00000000000000010010101001; 	// jal
disk[1385] <= 32'b000010_11110_11110_0000000000001000; 	// subi
disk[1386] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[1387] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1388] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[1389] <= 32'b111110_00000000000000001110010011; 	// jal
disk[1390] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1391] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[1392] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1393] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[1394] <= 32'b111100_00000000000000010101001100; 	// j
disk[1395] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[1396] <= 32'b010010_11101_10100_0000000001101010; 	// sw
disk[1397] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[1398] <= 32'b001110_11110_11100_0000000000000000; 	// mov
disk[1399] <= 32'b001110_11101_11011_0000000000000000; 	// mov
disk[1400] <= 32'b010000_00000_00000_0000000000000000; 	// li
disk[1401] <= 32'b010000_00000_11110_0000000000000000; 	// li
disk[1402] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[1403] <= 32'b000001_11110_11110_0000000111000000; 	// addi
disk[1404] <= 32'b010010_00000_00000_0000111111100000; 	// sw
disk[1405] <= 32'b010010_00000_00001_0000111111100001; 	// sw
disk[1406] <= 32'b010010_00000_00010_0000111111100010; 	// sw
disk[1407] <= 32'b010010_00000_00011_0000111111100011; 	// sw
disk[1408] <= 32'b010010_00000_00100_0000111111100100; 	// sw
disk[1409] <= 32'b010010_00000_00101_0000111111100101; 	// sw
disk[1410] <= 32'b010010_00000_00110_0000111111100110; 	// sw
disk[1411] <= 32'b010010_00000_00111_0000111111100111; 	// sw
disk[1412] <= 32'b010010_00000_01000_0000111111101000; 	// sw
disk[1413] <= 32'b010010_00000_01001_0000111111101001; 	// sw
disk[1414] <= 32'b010010_00000_01010_0000111111101010; 	// sw
disk[1415] <= 32'b010010_00000_01011_0000111111101011; 	// sw
disk[1416] <= 32'b010010_00000_01100_0000111111101100; 	// sw
disk[1417] <= 32'b010010_00000_01101_0000111111101101; 	// sw
disk[1418] <= 32'b010010_00000_01110_0000111111101110; 	// sw
disk[1419] <= 32'b010010_00000_01111_0000111111101111; 	// sw
disk[1420] <= 32'b010010_00000_10000_0000111111110000; 	// sw
disk[1421] <= 32'b010010_00000_10001_0000111111110001; 	// sw
disk[1422] <= 32'b010010_00000_10010_0000111111110010; 	// sw
disk[1423] <= 32'b010010_00000_10011_0000111111110011; 	// sw
disk[1424] <= 32'b010010_00000_10100_0000111111110100; 	// sw
disk[1425] <= 32'b010010_00000_10101_0000111111110101; 	// sw
disk[1426] <= 32'b010010_00000_10110_0000111111110110; 	// sw
disk[1427] <= 32'b010010_00000_10111_0000111111110111; 	// sw
disk[1428] <= 32'b010010_00000_11000_0000111111111000; 	// sw
disk[1429] <= 32'b010010_00000_11111_0000111111111001; 	// sw
disk[1430] <= 32'b001111_11110_00101_1111111111111011; 	// lw
disk[1431] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[1432] <= 32'b000000_00101_10000_01111_00000_001100; 	// eq
disk[1433] <= 32'b010101_01111_00000_0000010110100011; 	// jf
disk[1434] <= 32'b111110_00000000000000001001011001; 	// jal
disk[1435] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[1436] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1437] <= 32'b001111_11101_00110_0000000110101011; 	// lw
disk[1438] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1439] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[1440] <= 32'b010000_00000_10001_0000000000000001; 	// li
disk[1441] <= 32'b010010_11110_10001_1111111111111011; 	// sw
disk[1442] <= 32'b100110_00000_00000_0000000000000000; 	// cic
disk[1443] <= 32'b100101_00000_10010_0000000000000000; 	// gic
disk[1444] <= 32'b010010_11110_10010_1111111111111010; 	// sw
disk[1445] <= 32'b001111_11110_00101_1111111111111010; 	// lw
disk[1446] <= 32'b001111_11101_00110_0000000101110101; 	// lw
disk[1447] <= 32'b000000_00101_00110_10011_00000_001100; 	// eq
disk[1448] <= 32'b010101_10011_00000_0000011000100000; 	// jf
disk[1449] <= 32'b001110_11100_10100_0000000000000000; 	// mov
disk[1450] <= 32'b010010_11101_10100_0000000011110011; 	// sw
disk[1451] <= 32'b001111_11101_00111_0000000011110011; 	// lw
disk[1452] <= 32'b001111_11101_01000_0000000011110010; 	// lw
disk[1453] <= 32'b000000_00111_01000_10101_00000_000001; 	// sub
disk[1454] <= 32'b000001_10101_10110_0000000000000001; 	// addi
disk[1455] <= 32'b010010_11110_10110_0000000000000000; 	// sw
disk[1456] <= 32'b010001_11101_01001_0000000000011000; 	// la
disk[1457] <= 32'b001111_11101_01010_0000000001011111; 	// lw
disk[1458] <= 32'b000000_01001_01010_10111_00000_000000; 	// add
disk[1459] <= 32'b001111_11110_01011_0000000000000000; 	// lw
disk[1460] <= 32'b010010_10111_01011_0000000000000000; 	// sw
disk[1461] <= 32'b010001_11101_01100_0000000000000100; 	// la
disk[1462] <= 32'b000000_01100_01010_01111_00000_000000; 	// add
disk[1463] <= 32'b001111_11101_01101_0000000000000010; 	// lw
disk[1464] <= 32'b010010_01111_01101_0000000000000000; 	// sw
disk[1465] <= 32'b100111_00000_10000_0000000000000000; 	// gip
disk[1466] <= 32'b010001_11101_01110_0000000000001110; 	// la
disk[1467] <= 32'b000000_01110_01010_10001_00000_000000; 	// add
disk[1468] <= 32'b010010_10001_10000_0000000000000000; 	// sw
disk[1469] <= 32'b010001_11101_00101_0000000001000000; 	// la
disk[1470] <= 32'b000000_00101_01010_10010_00000_000000; 	// add
disk[1471] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[1472] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[1473] <= 32'b000000_10010_10100_10011_00000_001100; 	// eq
disk[1474] <= 32'b010101_10011_00000_0000010111001101; 	// jf
disk[1475] <= 32'b111110_00000000000000001010111001; 	// jal
disk[1476] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[1477] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1478] <= 32'b010010_11110_00101_1111111111111100; 	// sw
disk[1479] <= 32'b010001_11101_00110_0000000001000000; 	// la
disk[1480] <= 32'b001111_11101_00111_0000000001011111; 	// lw
disk[1481] <= 32'b000000_00110_00111_10101_00000_000000; 	// add
disk[1482] <= 32'b001111_11110_01000_1111111111111100; 	// lw
disk[1483] <= 32'b010010_10101_01000_0000000000000000; 	// sw
disk[1484] <= 32'b111100_00000000000000010111010010; 	// j
disk[1485] <= 32'b010001_11101_00101_0000000001000000; 	// la
disk[1486] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[1487] <= 32'b000000_00101_00110_10110_00000_000000; 	// add
disk[1488] <= 32'b001111_10110_10110_0000000000000000; 	// lw
disk[1489] <= 32'b010010_11110_10110_1111111111111100; 	// sw
disk[1490] <= 32'b001111_11101_00101_0000000011110010; 	// lw
disk[1491] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[1492] <= 32'b001111_11110_00110_1111111111111100; 	// lw
disk[1493] <= 32'b001111_11101_00111_0000000011101011; 	// lw
disk[1494] <= 32'b000000_00110_00111_10111_00000_000010; 	// mul
disk[1495] <= 32'b010010_11110_10111_1111111111111111; 	// sw
disk[1496] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1497] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[1498] <= 32'b000000_00101_10000_01111_00000_010000; 	// gt
disk[1499] <= 32'b010101_01111_00000_0000010111101111; 	// jf
disk[1500] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[1501] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1502] <= 32'b001111_00001_10001_0000000000000000; 	// lw
disk[1503] <= 32'b010010_11110_10001_1111111111111101; 	// sw
disk[1504] <= 32'b001111_11110_00111_1111111111111101; 	// lw
disk[1505] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1506] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[1507] <= 32'b001110_01000_00010_0000000000000000; 	// mov
disk[1508] <= 32'b010010_00010_00001_0000000000000000; 	// sw
disk[1509] <= 32'b000001_00110_10010_0000000000000001; 	// addi
disk[1510] <= 32'b010010_11110_10010_1111111111111110; 	// sw
disk[1511] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[1512] <= 32'b000001_01000_10011_0000000000000001; 	// addi
disk[1513] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[1514] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[1515] <= 32'b000010_00101_10100_0000000000000001; 	// subi
disk[1516] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[1517] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1518] <= 32'b111100_00000000000000010111011000; 	// j
disk[1519] <= 32'b001111_11101_00101_0000000001011111; 	// lw
disk[1520] <= 32'b001111_11101_00110_0000000001011110; 	// lw
disk[1521] <= 32'b000000_00101_00110_10101_00000_001100; 	// eq
disk[1522] <= 32'b010101_10101_00000_0000010111111001; 	// jf
disk[1523] <= 32'b000001_00101_10110_0000000000000001; 	// addi
disk[1524] <= 32'b001110_10110_00001_0000000000000000; 	// mov
disk[1525] <= 32'b111110_00000000000000010010101001; 	// jal
disk[1526] <= 32'b000010_11110_11110_0000000000001000; 	// subi
disk[1527] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1528] <= 32'b111100_00000000000000011000010111; 	// j
disk[1529] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[1530] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1531] <= 32'b111110_00000000000000000001100011; 	// jal
disk[1532] <= 32'b000010_11110_11110_0000000000000110; 	// subi
disk[1533] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1534] <= 32'b010001_11101_00110_0000000000000100; 	// la
disk[1535] <= 32'b001111_11101_00111_0000000001011111; 	// lw
disk[1536] <= 32'b000000_00110_00111_10111_00000_000000; 	// add
disk[1537] <= 32'b001111_11101_01000_0000000000000010; 	// lw
disk[1538] <= 32'b010010_10111_01000_0000000000000000; 	// sw
disk[1539] <= 32'b000001_00111_01111_0000000000000001; 	// addi
disk[1540] <= 32'b001110_01111_00001_0000000000000000; 	// mov
disk[1541] <= 32'b111110_00000000000000001101001110; 	// jal
disk[1542] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[1543] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1544] <= 32'b001111_11101_00110_0000000001101010; 	// lw
disk[1545] <= 32'b010000_00000_10001_0000000000000001; 	// li
disk[1546] <= 32'b000000_00110_10001_10000_00000_001100; 	// eq
disk[1547] <= 32'b010101_10000_00000_0000011000010111; 	// jf
disk[1548] <= 32'b001111_11101_00111_0000000110101011; 	// lw
disk[1549] <= 32'b010010_11101_00111_0000000110110110; 	// sw
disk[1550] <= 32'b001111_11101_01000_0000000110110110; 	// lw
disk[1551] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[1552] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[1553] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[1554] <= 32'b010000_00000_11110_0000000111000000; 	// li
disk[1555] <= 32'b100110_00000_00000_0000000000000000; 	// cic
disk[1556] <= 32'b111110_00000000000000010101000000; 	// jal
disk[1557] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1558] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1559] <= 32'b001111_11101_00101_0000000110101011; 	// lw
disk[1560] <= 32'b010010_11101_00101_0000000110110110; 	// sw
disk[1561] <= 32'b001111_11101_00110_0000000110110110; 	// lw
disk[1562] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1563] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[1564] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[1565] <= 32'b010000_00000_11110_0000000111000000; 	// li
disk[1566] <= 32'b100110_00000_00000_0000000000000000; 	// cic
disk[1567] <= 32'b111100_00000000000000011010001100; 	// j
disk[1568] <= 32'b001111_11110_00101_1111111111111010; 	// lw
disk[1569] <= 32'b001111_11101_00110_0000000101110100; 	// lw
disk[1570] <= 32'b000000_00101_00110_10010_00000_001100; 	// eq
disk[1571] <= 32'b010101_10010_00000_0000011010001100; 	// jf
disk[1572] <= 32'b001110_11100_10011_0000000000000000; 	// mov
disk[1573] <= 32'b010010_11101_10011_0000000011110011; 	// sw
disk[1574] <= 32'b001111_11101_00111_0000000011110011; 	// lw
disk[1575] <= 32'b001111_11101_01000_0000000011110010; 	// lw
disk[1576] <= 32'b000000_00111_01000_10100_00000_000001; 	// sub
disk[1577] <= 32'b000001_10100_10101_0000000000000001; 	// addi
disk[1578] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[1579] <= 32'b010001_11101_01001_0000000000011000; 	// la
disk[1580] <= 32'b001111_11101_01010_0000000001011111; 	// lw
disk[1581] <= 32'b000000_01001_01010_10110_00000_000000; 	// add
disk[1582] <= 32'b001111_11110_01011_0000000000000000; 	// lw
disk[1583] <= 32'b010010_10110_01011_0000000000000000; 	// sw
disk[1584] <= 32'b010001_11101_01100_0000000000000100; 	// la
disk[1585] <= 32'b000000_01100_01010_10111_00000_000000; 	// add
disk[1586] <= 32'b001111_11101_01101_0000000000000010; 	// lw
disk[1587] <= 32'b010010_10111_01101_0000000000000000; 	// sw
disk[1588] <= 32'b100111_00000_01111_0000000000000000; 	// gip
disk[1589] <= 32'b010001_11101_01110_0000000000001110; 	// la
disk[1590] <= 32'b000000_01110_01010_10000_00000_000000; 	// add
disk[1591] <= 32'b010010_10000_01111_0000000000000000; 	// sw
disk[1592] <= 32'b010001_11101_00101_0000000001000000; 	// la
disk[1593] <= 32'b000000_00101_01010_10001_00000_000000; 	// add
disk[1594] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[1595] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[1596] <= 32'b000000_10001_10011_10010_00000_001100; 	// eq
disk[1597] <= 32'b010101_10010_00000_0000011001001000; 	// jf
disk[1598] <= 32'b111110_00000000000000001010111001; 	// jal
disk[1599] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[1600] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1601] <= 32'b010010_11110_00101_1111111111111100; 	// sw
disk[1602] <= 32'b010001_11101_00110_0000000001000000; 	// la
disk[1603] <= 32'b001111_11101_00111_0000000001011111; 	// lw
disk[1604] <= 32'b000000_00110_00111_10100_00000_000000; 	// add
disk[1605] <= 32'b001111_11110_01000_1111111111111100; 	// lw
disk[1606] <= 32'b010010_10100_01000_0000000000000000; 	// sw
disk[1607] <= 32'b111100_00000000000000011001001101; 	// j
disk[1608] <= 32'b010001_11101_00101_0000000001000000; 	// la
disk[1609] <= 32'b001111_11101_00110_0000000001011111; 	// lw
disk[1610] <= 32'b000000_00101_00110_10101_00000_000000; 	// add
disk[1611] <= 32'b001111_10101_10101_0000000000000000; 	// lw
disk[1612] <= 32'b010010_11110_10101_1111111111111100; 	// sw
disk[1613] <= 32'b001111_11101_00101_0000000011110010; 	// lw
disk[1614] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[1615] <= 32'b001111_11110_00110_1111111111111100; 	// lw
disk[1616] <= 32'b001111_11101_00111_0000000011101011; 	// lw
disk[1617] <= 32'b000000_00110_00111_10110_00000_000010; 	// mul
disk[1618] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[1619] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1620] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[1621] <= 32'b000000_00101_01111_10111_00000_010000; 	// gt
disk[1622] <= 32'b010101_10111_00000_0000011001101010; 	// jf
disk[1623] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[1624] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1625] <= 32'b001111_00001_10000_0000000000000000; 	// lw
disk[1626] <= 32'b010010_11110_10000_1111111111111101; 	// sw
disk[1627] <= 32'b001111_11110_00111_1111111111111101; 	// lw
disk[1628] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1629] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[1630] <= 32'b001110_01000_00010_0000000000000000; 	// mov
disk[1631] <= 32'b010010_00010_00001_0000000000000000; 	// sw
disk[1632] <= 32'b000001_00110_10001_0000000000000001; 	// addi
disk[1633] <= 32'b010010_11110_10001_1111111111111110; 	// sw
disk[1634] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[1635] <= 32'b000001_01000_10010_0000000000000001; 	// addi
disk[1636] <= 32'b010010_11110_10010_1111111111111111; 	// sw
disk[1637] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[1638] <= 32'b000010_00101_10011_0000000000000001; 	// subi
disk[1639] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[1640] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[1641] <= 32'b111100_00000000000000011001010011; 	// j
disk[1642] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[1643] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1644] <= 32'b111110_00000000000000000001100011; 	// jal
disk[1645] <= 32'b000010_11110_11110_0000000000000110; 	// subi
disk[1646] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1647] <= 32'b010001_11101_00110_0000000000000100; 	// la
disk[1648] <= 32'b001111_11101_00111_0000000001011111; 	// lw
disk[1649] <= 32'b000000_00110_00111_10100_00000_000000; 	// add
disk[1650] <= 32'b001111_11101_01000_0000000000000001; 	// lw
disk[1651] <= 32'b010010_10100_01000_0000000000000000; 	// sw
disk[1652] <= 32'b001111_11101_01001_0000000110101011; 	// lw
disk[1653] <= 32'b010010_11101_01001_0000000110110110; 	// sw
disk[1654] <= 32'b001111_11101_01010_0000000110110110; 	// lw
disk[1655] <= 32'b001110_01010_00001_0000000000000000; 	// mov
disk[1656] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[1657] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[1658] <= 32'b010000_00000_11110_0000000111000000; 	// li
disk[1659] <= 32'b100110_00000_00000_0000000000000000; 	// cic
disk[1660] <= 32'b000001_00111_10101_0000000000000001; 	// addi
disk[1661] <= 32'b001110_10101_00001_0000000000000000; 	// mov
disk[1662] <= 32'b111110_00000000000000001110100110; 	// jal
disk[1663] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1664] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1665] <= 32'b111110_00000000000000010101000000; 	// jal
disk[1666] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1667] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1668] <= 32'b001111_11101_00110_0000000110101011; 	// lw
disk[1669] <= 32'b010010_11101_00110_0000000110110110; 	// sw
disk[1670] <= 32'b001111_11101_00111_0000000110110110; 	// lw
disk[1671] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1672] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[1673] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[1674] <= 32'b010000_00000_11110_0000000111000000; 	// li
disk[1675] <= 32'b100110_00000_00000_0000000000000000; 	// cic
disk[1676] <= 32'b010000_00000_10110_0000000000000001; 	// li
disk[1677] <= 32'b010101_10110_00000_0000011110011000; 	// jf
disk[1678] <= 32'b010011_00000_10111_0000000000000000; 	// in
disk[1679] <= 32'b010010_11110_10111_1111111111111001; 	// sw
disk[1680] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1681] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1682] <= 32'b010000_00000_00010_0000000000000000; 	// li
disk[1683] <= 32'b010100_00000_00001_0000000000000000; 	// out
disk[1684] <= 32'b001111_11101_00110_0000000110110110; 	// lw
disk[1685] <= 32'b001111_11101_00111_0000000110101011; 	// lw
disk[1686] <= 32'b000000_00110_00111_01111_00000_001100; 	// eq
disk[1687] <= 32'b010101_01111_00000_0000011010111100; 	// jf
disk[1688] <= 32'b010000_00000_10001_0000000000000001; 	// li
disk[1689] <= 32'b000000_00101_10001_10000_00000_001100; 	// eq
disk[1690] <= 32'b010101_10000_00000_0000011010011111; 	// jf
disk[1691] <= 32'b001111_11101_01000_0000000110101100; 	// lw
disk[1692] <= 32'b010010_11110_01000_1111111111111001; 	// sw
disk[1693] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1694] <= 32'b111100_00000000000000011010111011; 	// j
disk[1695] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1696] <= 32'b010000_00000_10011_0000000000000010; 	// li
disk[1697] <= 32'b000000_00101_10011_10010_00000_001100; 	// eq
disk[1698] <= 32'b010101_10010_00000_0000011010100111; 	// jf
disk[1699] <= 32'b001111_11101_00110_0000000110101111; 	// lw
disk[1700] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1701] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1702] <= 32'b111100_00000000000000011010111011; 	// j
disk[1703] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1704] <= 32'b010000_00000_10101_0000000000000011; 	// li
disk[1705] <= 32'b000000_00101_10101_10100_00000_001100; 	// eq
disk[1706] <= 32'b010101_10100_00000_0000011010101111; 	// jf
disk[1707] <= 32'b001111_11101_00110_0000000110110010; 	// lw
disk[1708] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1709] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1710] <= 32'b111100_00000000000000011010111011; 	// j
disk[1711] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1712] <= 32'b010000_00000_10111_0000000000000100; 	// li
disk[1713] <= 32'b000000_00101_10111_10110_00000_001100; 	// eq
disk[1714] <= 32'b010101_10110_00000_0000011010111001; 	// jf
disk[1715] <= 32'b111110_00000000000000000000110011; 	// jal
disk[1716] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[1717] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1718] <= 32'b001111_11101_00110_0000000110101011; 	// lw
disk[1719] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1720] <= 32'b111100_00000000000000011010111011; 	// j
disk[1721] <= 32'b001111_11101_00101_0000000110101011; 	// lw
disk[1722] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1723] <= 32'b111100_00000000000000011110010010; 	// j
disk[1724] <= 32'b001111_11101_00101_0000000110110110; 	// lw
disk[1725] <= 32'b001111_11101_00110_0000000110101100; 	// lw
disk[1726] <= 32'b000000_00101_00110_01111_00000_001100; 	// eq
disk[1727] <= 32'b010101_01111_00000_0000011011100101; 	// jf
disk[1728] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1729] <= 32'b010000_00000_10001_0000000000000001; 	// li
disk[1730] <= 32'b000000_00111_10001_10000_00000_001100; 	// eq
disk[1731] <= 32'b010101_10000_00000_0000011011001000; 	// jf
disk[1732] <= 32'b001111_11101_01000_0000000110101011; 	// lw
disk[1733] <= 32'b010010_11110_01000_1111111111111001; 	// sw
disk[1734] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1735] <= 32'b111100_00000000000000011011100100; 	// j
disk[1736] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1737] <= 32'b010000_00000_10011_0000000000000010; 	// li
disk[1738] <= 32'b000000_00101_10011_10010_00000_001100; 	// eq
disk[1739] <= 32'b010101_10010_00000_0000011011010101; 	// jf
disk[1740] <= 32'b001111_11101_00110_0000000110101110; 	// lw
disk[1741] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1742] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1743] <= 32'b111110_00000000000000000100100000; 	// jal
disk[1744] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1745] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1746] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1747] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[1748] <= 32'b111100_00000000000000011011100100; 	// j
disk[1749] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1750] <= 32'b010000_00000_10101_0000000000000011; 	// li
disk[1751] <= 32'b000000_00101_10101_10100_00000_001100; 	// eq
disk[1752] <= 32'b010101_10100_00000_0000011011100010; 	// jf
disk[1753] <= 32'b001111_11101_00110_0000000110101101; 	// lw
disk[1754] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1755] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1756] <= 32'b111110_00000000000000000100100000; 	// jal
disk[1757] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1758] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1759] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1760] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[1761] <= 32'b111100_00000000000000011011100100; 	// j
disk[1762] <= 32'b001111_11101_00101_0000000110101011; 	// lw
disk[1763] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1764] <= 32'b111100_00000000000000011110010010; 	// j
disk[1765] <= 32'b001111_11101_00101_0000000110110110; 	// lw
disk[1766] <= 32'b001111_11101_00110_0000000110101101; 	// lw
disk[1767] <= 32'b000000_00101_00110_10110_00000_001100; 	// eq
disk[1768] <= 32'b010101_10110_00000_0000011011110100; 	// jf
disk[1769] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1770] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[1771] <= 32'b000000_00111_01111_10111_00000_010000; 	// gt
disk[1772] <= 32'b010101_10111_00000_0000011011110001; 	// jf
disk[1773] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1774] <= 32'b111110_00000000000000000011001111; 	// jal
disk[1775] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[1776] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1777] <= 32'b001111_11101_00101_0000000110101011; 	// lw
disk[1778] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1779] <= 32'b111100_00000000000000011110010010; 	// j
disk[1780] <= 32'b001111_11101_00101_0000000110110110; 	// lw
disk[1781] <= 32'b001111_11101_00110_0000000110101110; 	// lw
disk[1782] <= 32'b000000_00101_00110_10000_00000_001100; 	// eq
disk[1783] <= 32'b010101_10000_00000_0000011100000011; 	// jf
disk[1784] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1785] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[1786] <= 32'b000000_00111_10010_10001_00000_010000; 	// gt
disk[1787] <= 32'b010101_10001_00000_0000011100000000; 	// jf
disk[1788] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1789] <= 32'b111110_00000000000000000100001110; 	// jal
disk[1790] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1791] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1792] <= 32'b001111_11101_00101_0000000110101011; 	// lw
disk[1793] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1794] <= 32'b111100_00000000000000011110010010; 	// j
disk[1795] <= 32'b001111_11101_00101_0000000110110110; 	// lw
disk[1796] <= 32'b001111_11101_00110_0000000110101111; 	// lw
disk[1797] <= 32'b000000_00101_00110_10011_00000_001100; 	// eq
disk[1798] <= 32'b010101_10011_00000_0000011100101100; 	// jf
disk[1799] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1800] <= 32'b010000_00000_10101_0000000000000001; 	// li
disk[1801] <= 32'b000000_00111_10101_10100_00000_001100; 	// eq
disk[1802] <= 32'b010101_10100_00000_0000011100010100; 	// jf
disk[1803] <= 32'b001111_11101_01000_0000000110110000; 	// lw
disk[1804] <= 32'b010010_11110_01000_1111111111111001; 	// sw
disk[1805] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1806] <= 32'b111110_00000000000000000100100000; 	// jal
disk[1807] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1808] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1809] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1810] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[1811] <= 32'b111100_00000000000000011100101011; 	// j
disk[1812] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1813] <= 32'b010000_00000_10111_0000000000000010; 	// li
disk[1814] <= 32'b000000_00101_10111_10110_00000_001100; 	// eq
disk[1815] <= 32'b010101_10110_00000_0000011100011100; 	// jf
disk[1816] <= 32'b001111_11101_00110_0000000110101011; 	// lw
disk[1817] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1818] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1819] <= 32'b111100_00000000000000011100101011; 	// j
disk[1820] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1821] <= 32'b010000_00000_10000_0000000000000011; 	// li
disk[1822] <= 32'b000000_00101_10000_01111_00000_001100; 	// eq
disk[1823] <= 32'b010101_01111_00000_0000011100101001; 	// jf
disk[1824] <= 32'b001111_11101_00110_0000000110110001; 	// lw
disk[1825] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1826] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1827] <= 32'b111110_00000000000000001011110101; 	// jal
disk[1828] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1829] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1830] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1831] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[1832] <= 32'b111100_00000000000000011100101011; 	// j
disk[1833] <= 32'b001111_11101_00101_0000000110101011; 	// lw
disk[1834] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1835] <= 32'b111100_00000000000000011110010010; 	// j
disk[1836] <= 32'b001111_11101_00101_0000000110110110; 	// lw
disk[1837] <= 32'b001111_11101_00110_0000000110110000; 	// lw
disk[1838] <= 32'b000000_00101_00110_10001_00000_001100; 	// eq
disk[1839] <= 32'b010101_10001_00000_0000011100111011; 	// jf
disk[1840] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1841] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[1842] <= 32'b000000_00111_10011_10010_00000_010000; 	// gt
disk[1843] <= 32'b010101_10010_00000_0000011100111000; 	// jf
disk[1844] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1845] <= 32'b111110_00000000000000010000010110; 	// jal
disk[1846] <= 32'b000010_11110_11110_0000000000001010; 	// subi
disk[1847] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1848] <= 32'b001111_11101_00101_0000000110101011; 	// lw
disk[1849] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1850] <= 32'b111100_00000000000000011110010010; 	// j
disk[1851] <= 32'b001111_11101_00101_0000000110110110; 	// lw
disk[1852] <= 32'b001111_11101_00110_0000000110110001; 	// lw
disk[1853] <= 32'b000000_00101_00110_10100_00000_001100; 	// eq
disk[1854] <= 32'b010101_10100_00000_0000011101001010; 	// jf
disk[1855] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1856] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[1857] <= 32'b000000_00111_10110_10101_00000_010000; 	// gt
disk[1858] <= 32'b010101_10101_00000_0000011101000111; 	// jf
disk[1859] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1860] <= 32'b111110_00000000000000000010000110; 	// jal
disk[1861] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[1862] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1863] <= 32'b001111_11101_00101_0000000110101011; 	// lw
disk[1864] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1865] <= 32'b111100_00000000000000011110010010; 	// j
disk[1866] <= 32'b001111_11101_00101_0000000110110110; 	// lw
disk[1867] <= 32'b001111_11101_00110_0000000110110010; 	// lw
disk[1868] <= 32'b000000_00101_00110_10111_00000_001100; 	// eq
disk[1869] <= 32'b010101_10111_00000_0000011101110101; 	// jf
disk[1870] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1871] <= 32'b010000_00000_10000_0000000000000001; 	// li
disk[1872] <= 32'b000000_00111_10000_01111_00000_001100; 	// eq
disk[1873] <= 32'b010101_01111_00000_0000011101011010; 	// jf
disk[1874] <= 32'b010000_00000_10001_0000000000000001; 	// li
disk[1875] <= 32'b010010_11101_10001_0000000001101010; 	// sw
disk[1876] <= 32'b111110_00000000000000010101000000; 	// jal
disk[1877] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1878] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1879] <= 32'b001111_11101_00110_0000000110101011; 	// lw
disk[1880] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1881] <= 32'b111100_00000000000000011101110100; 	// j
disk[1882] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1883] <= 32'b010000_00000_10011_0000000000000010; 	// li
disk[1884] <= 32'b000000_00101_10011_10010_00000_001100; 	// eq
disk[1885] <= 32'b010101_10010_00000_0000011101100110; 	// jf
disk[1886] <= 32'b111110_00000000000000001011110101; 	// jal
disk[1887] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1888] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1889] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1890] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[1891] <= 32'b001111_11101_00110_0000000110110011; 	// lw
disk[1892] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1893] <= 32'b111100_00000000000000011101110100; 	// j
disk[1894] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1895] <= 32'b010000_00000_10101_0000000000000011; 	// li
disk[1896] <= 32'b000000_00101_10101_10100_00000_001100; 	// eq
disk[1897] <= 32'b010101_10100_00000_0000011101110010; 	// jf
disk[1898] <= 32'b111110_00000000000000001100010110; 	// jal
disk[1899] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[1900] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1901] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[1902] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[1903] <= 32'b001111_11101_00110_0000000110110100; 	// lw
disk[1904] <= 32'b010010_11110_00110_1111111111111001; 	// sw
disk[1905] <= 32'b111100_00000000000000011101110100; 	// j
disk[1906] <= 32'b001111_11101_00101_0000000110101011; 	// lw
disk[1907] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1908] <= 32'b111100_00000000000000011110010010; 	// j
disk[1909] <= 32'b001111_11101_00101_0000000110110110; 	// lw
disk[1910] <= 32'b001111_11101_00110_0000000110110011; 	// lw
disk[1911] <= 32'b000000_00101_00110_10110_00000_001100; 	// eq
disk[1912] <= 32'b010101_10110_00000_0000011110000100; 	// jf
disk[1913] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1914] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[1915] <= 32'b000000_00111_01111_10111_00000_010000; 	// gt
disk[1916] <= 32'b010101_10111_00000_0000011110000001; 	// jf
disk[1917] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1918] <= 32'b111110_00000000000000010100110010; 	// jal
disk[1919] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1920] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1921] <= 32'b001111_11101_00101_0000000110101011; 	// lw
disk[1922] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1923] <= 32'b111100_00000000000000011110010010; 	// j
disk[1924] <= 32'b001111_11101_00101_0000000110110110; 	// lw
disk[1925] <= 32'b001111_11101_00110_0000000110110100; 	// lw
disk[1926] <= 32'b000000_00101_00110_10000_00000_001100; 	// eq
disk[1927] <= 32'b010101_10000_00000_0000011110010010; 	// jf
disk[1928] <= 32'b001111_11110_00111_1111111111111001; 	// lw
disk[1929] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[1930] <= 32'b000000_00111_10010_10001_00000_010000; 	// gt
disk[1931] <= 32'b010101_10001_00000_0000011110010000; 	// jf
disk[1932] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[1933] <= 32'b111110_00000000000000010100011110; 	// jal
disk[1934] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[1935] <= 32'b001110_11000_00101_0000000000000000; 	// mov
disk[1936] <= 32'b001111_11101_00101_0000000110101011; 	// lw
disk[1937] <= 32'b010010_11110_00101_1111111111111001; 	// sw
disk[1938] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[1939] <= 32'b010010_11101_00101_0000000110110110; 	// sw
disk[1940] <= 32'b001111_11101_00110_0000000110110110; 	// lw
disk[1941] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[1942] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[1943] <= 32'b111100_00000000000000011010001100; 	// j
disk[1944] <= 32'b111111_00000000000000000000000000; 	// halt


		// PROGRAMA 1
		disk[3800] <= 32'b111101_00000000000000000000100011;		// Jump to Main
		disk[3801] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[3802] <= 32'b010010_11110_00001_1111111111111100; 	// sw
		disk[3803] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[3804] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[3805] <= 32'b010000_00000_10000_0000000000000001; 	// li
		disk[3806] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[3807] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[3808] <= 32'b010010_11110_10001_1111111111111101; 	// sw
		disk[3809] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[3810] <= 32'b001111_11110_00110_1111111111111100; 	// lw
		disk[3811] <= 32'b000000_00101_00110_10010_00000_001111; 	// let
		disk[3812] <= 32'b010101_10010_00000_0000000000100000; 	// jf
		disk[3813] <= 32'b010000_00000_10100_0000000000000001; 	// li
		disk[3814] <= 32'b000000_00101_10100_10011_00000_001111; 	// let
		disk[3815] <= 32'b010101_10011_00000_0000000000010010; 	// jf
		disk[3816] <= 32'b010010_11110_00101_1111111111111110; 	// sw
		disk[3817] <= 32'b111100_00000000000000000000011011; 	// j
		disk[3818] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[3819] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[3820] <= 32'b000000_00101_00110_10101_00000_000000; 	// add
		disk[3821] <= 32'b010010_11110_10101_1111111111111110; 	// sw
		disk[3822] <= 32'b010010_11110_00110_1111111111111111; 	// sw
		disk[3823] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[3824] <= 32'b001111_11110_00111_1111111111111110; 	// lw
		disk[3825] <= 32'b010010_11110_00111_0000000000000000; 	// sw
		disk[3826] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[3827] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[3828] <= 32'b000001_00101_10110_0000000000000001; 	// addi
		disk[3829] <= 32'b010010_11110_10110_1111111111111101; 	// sw
		disk[3830] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[3831] <= 32'b111100_00000000000000000000001001; 	// j
		disk[3832] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[3833] <= 32'b001110_00101_11000_0000000000000000; 	// mov
		disk[3834] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[3835] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[3836] <= 32'b010000_00000_01111_0000000000001011; 	// li
		disk[3837] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[3838] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[3839] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[3840] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[3841] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[3842] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[3843] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[3844] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[3845] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[3846] <= 32'b010000_00000_00010_0000000000000000; 	// li
		disk[3847] <= 32'b010100_00000_00001_0000000000000000; 	// out
		disk[3848] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[3849] <= 32'b011111_11001_00000_0000000000000000; 	// syscall
		
		// PROGRAMA 2
		disk[3900] <= 32'b111101_00000000000000000000100001;		// Jump to Main
		disk[3901] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[3902] <= 32'b010010_11110_00001_1111111111111100; 	// sw
		disk[3903] <= 32'b010010_11110_00010_1111111111111101; 	// sw
		disk[3904] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[3905] <= 32'b010010_11110_01111_1111111111111110; 	// sw
		disk[3906] <= 32'b010000_00000_10000_0000000000000000; 	// li
		disk[3907] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[3908] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[3909] <= 32'b001111_11110_00110_1111111111111101; 	// lw
		disk[3910] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
		disk[3911] <= 32'b010101_10001_00000_0000000000011100; 	// jf
		disk[3912] <= 32'b001111_11110_00111_1111111111111100; 	// lw
		disk[3913] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
		disk[3914] <= 32'b001111_10010_10010_0000000000000000; 	// lw
		disk[3915] <= 32'b001111_11110_01000_0000000000000000; 	// lw
		disk[3916] <= 32'b000000_01000_10010_10011_00000_001110; 	// lt
		disk[3917] <= 32'b010101_10011_00000_0000000000010111; 	// jf
		disk[3918] <= 32'b000000_00111_00101_10100_00000_000000; 	// add
		disk[3919] <= 32'b001111_10100_10100_0000000000000000; 	// lw
		disk[3920] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[3921] <= 32'b001111_11110_01000_0000000000000000; 	// lw
		disk[3922] <= 32'b010010_11110_00101_1111111111111111; 	// sw
		disk[3923] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[3924] <= 32'b000001_00101_10101_0000000000000001; 	// addi
		disk[3925] <= 32'b010010_11110_10101_1111111111111110; 	// sw
		disk[3926] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[3927] <= 32'b111100_00000000000000000000001000; 	// j
		disk[3928] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[3929] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[3930] <= 32'b010000_00000_00010_0000000000000001; 	// li
		disk[3931] <= 32'b010100_00000_00001_0000000000000001; 	// out
		disk[3932] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[3933] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[3934] <= 32'b010001_11110_00101_1111111111111011; 	// la
		disk[3935] <= 32'b010000_00000_01111_0000000000001100; 	// li
		disk[3936] <= 32'b010010_00101_01111_0000000000000000; 	// sw
		disk[3937] <= 32'b010000_00000_10000_0000000000101001; 	// li
		disk[3938] <= 32'b010010_00101_10000_0000000000000001; 	// sw
		disk[3939] <= 32'b010000_00000_10001_0000000000010111; 	// li
		disk[3940] <= 32'b010010_00101_10001_0000000000000010; 	// sw
		disk[3941] <= 32'b010000_00000_10010_0000000001100010; 	// li
		disk[3942] <= 32'b010010_00101_10010_0000000000000011; 	// sw
		disk[3943] <= 32'b010000_00000_10011_0000000000100001; 	// li
		disk[3944] <= 32'b010010_00101_10011_0000000000000100; 	// sw
		disk[3945] <= 32'b010000_00000_10100_0000000000010101; 	// li
		disk[3946] <= 32'b010010_00101_10100_0000000000000101; 	// sw
		disk[3947] <= 32'b010001_11110_00001_1111111111111011; 	// la
		disk[3948] <= 32'b010000_00000_00010_0000000000000110; 	// li
		disk[3949] <= 32'b010010_11110_11111_1111111111111010; 	// sw
		disk[3950] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[3951] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[3952] <= 32'b001111_11110_11111_1111111111111010; 	// lw
		disk[3953] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[3954] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[3955] <= 32'b011111_11001_00000_0000000000000000; 	// syscall
		
		// PROGRAMA 3
		disk[4000] <= 32'b111101_00000000000000000000010100;		// Jump to Main
		disk[4001] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[4002] <= 32'b010010_11110_00001_1111111111111111; 	// sw
		disk[4003] <= 32'b010000_00000_01111_0000000000000001; 	// li
		disk[4004] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[4005] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[4006] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[4007] <= 32'b000000_00101_10001_10000_00000_010000; 	// gt
		disk[4008] <= 32'b010101_10000_00000_0000000000010001; 	// jf
		disk[4009] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[4010] <= 32'b000000_00110_00101_10010_00000_000010; 	// mul
		disk[4011] <= 32'b010010_11110_10010_0000000000000000; 	// sw
		disk[4012] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[4013] <= 32'b000010_00101_10011_0000000000000001; 	// subi
		disk[4014] <= 32'b010010_11110_10011_1111111111111111; 	// sw
		disk[4015] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[4016] <= 32'b111100_00000000000000000000000101; 	// j
		disk[4017] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[4018] <= 32'b001110_00101_11000_0000000000000000; 	// mov
		disk[4019] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[4020] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[4021] <= 32'b010000_00000_01111_0000000001011101; 	// li
		disk[4022] <= 32'b010010_11110_01111_1111111111111110; 	// sw
		disk[4023] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[4024] <= 32'b010010_11110_00101_1111111111111111; 	// sw
		disk[4025] <= 32'b101000_00000000000000000000000000; 	// preIO
		disk[4026] <= 32'b010011_00000_10000_0000000000000000; 	// in
		disk[4027] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[4028] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[4029] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[4030] <= 32'b010010_11110_11111_1111111111111101; 	// sw
		disk[4031] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[4032] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[4033] <= 32'b001111_11110_11111_1111111111111101; 	// lw
		disk[4034] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[4035] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[4036] <= 32'b010000_00000_00010_0000000000000010; 	// li
		disk[4037] <= 32'b010100_00000_00001_0000000000000010; 	// out
		disk[4038] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[4039] <= 32'b011111_11001_00000_0000000000000000; 	// syscall
		
	end
endmodule
