module disco_rigido (clk, we, addr, datain, dataout);
	input clk;										// clock
	input we;										// write enable
	input [31:0] addr;							// disk address
	input [31:0] datain;							// data in (to disk)
	
	output reg [31:0] dataout;					// data out (from disk)
	
	localparam DISK_SIZE = 500;				// Tamanho do disco
	reg [31:0] disk [DISK_SIZE-1:0];			// disk cells
	
	always @ (posedge clk) begin
		if (we) disk[addr] <= datain;			// write disk
	end
	
	always @ (negedge clk) begin
		dataout <= disk[addr];
	end

	initial begin
		// SISTEMA OPERACIONAL
disk[0] <= 32'b010110_00000000000000000010000100;		// Jump to Main
disk[1] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[2] <= 32'b010000_00000_10100_0000000000100000; 	// li
disk[3] <= 32'b010010_00101_10100_0000000000100000; 	// sw
disk[4] <= 32'b010000_00000_10101_0000000001100100; 	// li
disk[5] <= 32'b010010_00101_10101_0000000000100001; 	// sw
disk[6] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[7] <= 32'b010010_11110_10110_0000000000000000; 	// sw
disk[8] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[9] <= 32'b010000_00000_11000_0000000000100000; 	// li
disk[10] <= 32'b000000_01010_11000_10111_00000_001110; 	// lt
disk[11] <= 32'b010101_10111_00000_0000000000010100; 	// jf
disk[12] <= 32'b010001_00101_01011_0000000000000000; 	// la
disk[13] <= 32'b000000_01011_01010_11001_00000_000000; 	// add
disk[14] <= 32'b010000_00000_11010_0000000000000000; 	// li
disk[15] <= 32'b010010_11001_11010_0000000000000000; 	// sw
disk[16] <= 32'b000001_01010_11011_0000000000000001; 	// addi
disk[17] <= 32'b010010_11110_11011_0000000000000000; 	// sw
disk[18] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[19] <= 32'b010110_00000000000000000000001000; 	// j
disk[20] <= 32'b010000_00000_11100_0000000000000000; 	// li
disk[21] <= 32'b010010_11110_11100_0000000000000000; 	// sw
disk[22] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[23] <= 32'b010000_00000_10100_0000000000000111; 	// li
disk[24] <= 32'b000000_01010_10100_11101_00000_001110; 	// lt
disk[25] <= 32'b010101_11101_00000_0000000000100001; 	// jf
disk[26] <= 32'b000000_01011_01010_10101_00000_000000; 	// add
disk[27] <= 32'b010000_00000_10110_0000000000000001; 	// li
disk[28] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[29] <= 32'b000001_01010_10111_0000000000000001; 	// addi
disk[30] <= 32'b010010_11110_10111_0000000000000000; 	// sw
disk[31] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[32] <= 32'b010110_00000000000000000000010111; 	// j
disk[33] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[34] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[35] <= 32'b010000_00000_00110_0000000000000000; 	// li
disk[36] <= 32'b010000_00000_00111_0000000000000000; 	// li
disk[37] <= 32'b010100_00000_00110_0000000000000000; 	// out
disk[38] <= 32'b010000_00000_00110_0000000000000000; 	// li
disk[39] <= 32'b010000_00000_00111_0000000000000001; 	// li
disk[40] <= 32'b010100_00000_00110_0000000000000001; 	// out
disk[41] <= 32'b010000_00000_00110_0000000000000000; 	// li
disk[42] <= 32'b010000_00000_00111_0000000000000010; 	// li
disk[43] <= 32'b010100_00000_00110_0000000000000010; 	// out
disk[44] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[45] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[46] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[47] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[48] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[49] <= 32'b010000_00000_10110_0000000000100000; 	// li
disk[50] <= 32'b000000_01010_10110_10101_00000_001110; 	// lt
disk[51] <= 32'b010101_10101_00000_0000000001001011; 	// jf
disk[52] <= 32'b010001_00101_01011_0000000000000000; 	// la
disk[53] <= 32'b000000_01011_01010_10111_00000_000000; 	// add
disk[54] <= 32'b001111_10111_10111_0000000000000000; 	// lw
disk[55] <= 32'b010000_00000_11001_0000000000000000; 	// li
disk[56] <= 32'b000000_10111_11001_11000_00000_001100; 	// eq
disk[57] <= 32'b010101_11000_00000_0000000001000111; 	// jf
disk[58] <= 32'b000000_01011_01010_11010_00000_000000; 	// add
disk[59] <= 32'b010000_00000_11011_0000000000000001; 	// li
disk[60] <= 32'b010010_11010_11011_0000000000000000; 	// sw
disk[61] <= 32'b000001_01010_11100_0000000000000001; 	// addi
disk[62] <= 32'b000000_01011_11100_11101_00000_000000; 	// add
disk[63] <= 32'b010000_00000_10100_0000000000000001; 	// li
disk[64] <= 32'b010010_11101_10100_0000000000000000; 	// sw
disk[65] <= 32'b000001_01010_10101_0000000000000010; 	// addi
disk[66] <= 32'b000000_01011_10101_10110_00000_000000; 	// add
disk[67] <= 32'b010000_00000_10111_0000000000000001; 	// li
disk[68] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[69] <= 32'b001110_01010_00001_0000000000000000; 	// mov
disk[70] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[71] <= 32'b000001_01010_11000_0000000000000001; 	// addi
disk[72] <= 32'b010010_11110_11000_0000000000000000; 	// sw
disk[73] <= 32'b001111_11110_01010_0000000000000000; 	// lw
disk[74] <= 32'b010110_00000000000000000000110000; 	// j
disk[75] <= 32'b001111_00101_01100_0000000000100001; 	// lw
disk[76] <= 32'b001110_01100_00001_0000000000000000; 	// mov
disk[77] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[78] <= 32'b000001_11110_11110_0000000000001001; 	// addi
disk[79] <= 32'b010010_11110_00110_1111111111111010; 	// sw
disk[80] <= 32'b010010_11110_00111_1111111111111011; 	// sw
disk[81] <= 32'b010000_00000_10100_0000000000100101; 	// li
disk[82] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[83] <= 32'b001111_11110_01010_1111111111111010; 	// lw
disk[84] <= 32'b010010_11110_01010_1111111111111100; 	// sw
disk[85] <= 32'b010010_11110_01010_1111111111111010; 	// sw
disk[86] <= 32'b010010_11110_11111_1111111111111001; 	// sw
disk[87] <= 32'b010111_00000000000000000000101101; 	// jal
disk[88] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[89] <= 32'b001111_11110_01010_1111111111111010; 	// lw
disk[90] <= 32'b001111_11110_11111_1111111111111001; 	// lw
disk[91] <= 32'b001110_00001_01011_0000000000000000; 	// mov
disk[92] <= 32'b010010_11110_01011_1111111111111111; 	// sw
disk[93] <= 32'b001111_00101_01100_0000000000100000; 	// lw
disk[94] <= 32'b001111_11110_01101_1111111111111111; 	// lw
disk[95] <= 32'b000000_01100_01101_10101_00000_000010; 	// mul
disk[96] <= 32'b010010_11110_10101_1111111111111101; 	// sw
disk[97] <= 32'b001111_11110_01110_1111111111111100; 	// lw
disk[98] <= 32'b001110_01110_00110_0000000000000000; 	// mov
disk[99] <= 32'b011001_00110_10110_0000000000000000; 	// ldk
disk[100] <= 32'b010010_11110_10110_1111111111111110; 	// sw
disk[101] <= 32'b001111_11110_01111_1111111111111110; 	// lw
disk[102] <= 32'b001101_01111_10111_0000000000011010; 	// srli
disk[103] <= 32'b001111_11110_10000_0000000000000000; 	// lw
disk[104] <= 32'b000000_10111_10000_11000_00000_001101; 	// ne
disk[105] <= 32'b010101_11000_00000_0000000001111001; 	// jf
disk[106] <= 32'b001110_01111_00110_0000000000000000; 	// mov
disk[107] <= 32'b001111_11110_10001_1111111111111101; 	// lw
disk[108] <= 32'b001110_10001_00111_0000000000000000; 	// mov
disk[109] <= 32'b011100_00111_00110_0000000000000000; 	// sim
disk[110] <= 32'b000001_01110_11001_0000000000000001; 	// addi
disk[111] <= 32'b010010_11110_11001_1111111111111100; 	// sw
disk[112] <= 32'b001111_11110_01110_1111111111111100; 	// lw
disk[113] <= 32'b001110_01110_00110_0000000000000000; 	// mov
disk[114] <= 32'b011001_00110_11010_0000000000000000; 	// ldk
disk[115] <= 32'b010010_11110_11010_1111111111111110; 	// sw
disk[116] <= 32'b001111_11110_01111_1111111111111110; 	// lw
disk[117] <= 32'b000001_10001_11011_0000000000000001; 	// addi
disk[118] <= 32'b010010_11110_11011_1111111111111101; 	// sw
disk[119] <= 32'b001111_11110_10001_1111111111111101; 	// lw
disk[120] <= 32'b010110_00000000000000000001100101; 	// j
disk[121] <= 32'b001110_01111_00110_0000000000000000; 	// mov
disk[122] <= 32'b001110_10001_00111_0000000000000000; 	// mov
disk[123] <= 32'b011100_00111_00110_0000000000000000; 	// sim
disk[124] <= 32'b001111_11110_10010_1111111111111011; 	// lw
disk[125] <= 32'b001110_10010_00110_0000000000000000; 	// mov
disk[126] <= 32'b100100_00110_00000_0000000000000000; 	// mmuSelect
disk[127] <= 32'b000000_01100_01101_11100_00000_000010; 	// mul
disk[128] <= 32'b001110_11100_00110_0000000000000000; 	// mov
disk[129] <= 32'b100000_00000_00110_0000000000000000; 	// mmuLowerIM
disk[130] <= 32'b001110_10001_00001_0000000000000000; 	// mov
disk[131] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[132] <= 32'b001110_00000_00101_0000000000000000; 	// mov
disk[133] <= 32'b000001_11110_11110_0000000000100110; 	// addi
disk[134] <= 32'b010010_11110_11111_1111111111111101; 	// sw
disk[135] <= 32'b010111_00000000000000000000000001; 	// jal
disk[136] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[137] <= 32'b001111_11110_11111_1111111111111101; 	// lw
disk[138] <= 32'b001110_00001_01010_0000000000000000; 	// mov
disk[139] <= 32'b010000_00000_10100_0000000011111010; 	// li
disk[140] <= 32'b010010_11110_10100_1111111111111110; 	// sw
disk[141] <= 32'b010000_00000_10101_0000000100101100; 	// li
disk[142] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[143] <= 32'b010000_00000_10110_0000000101100010; 	// li
disk[144] <= 32'b010010_11110_10110_0000000000000000; 	// sw
disk[145] <= 32'b001111_11110_01011_1111111111111110; 	// lw
disk[146] <= 32'b001110_01011_00110_0000000000000000; 	// mov
disk[147] <= 32'b010000_00000_00111_0000000000000001; 	// li
disk[148] <= 32'b010010_11110_01010_1111111111111001; 	// sw
disk[149] <= 32'b010010_11110_11111_1111111111111101; 	// sw
disk[150] <= 32'b010111_00000000000000000001001110; 	// jal
disk[151] <= 32'b000010_11110_11110_0000000000001001; 	// subi
disk[152] <= 32'b001111_11110_01010_1111111111111001; 	// lw
disk[153] <= 32'b001111_11110_11111_1111111111111101; 	// lw
disk[154] <= 32'b001110_00001_01100_0000000000000000; 	// mov
disk[155] <= 32'b001111_11110_01101_1111111111111111; 	// lw
disk[156] <= 32'b001110_01101_00110_0000000000000000; 	// mov
disk[157] <= 32'b010000_00000_00111_0000000000000010; 	// li
disk[158] <= 32'b010010_11110_01010_1111111111111001; 	// sw
disk[159] <= 32'b010010_11110_01100_1111111111111001; 	// sw
disk[160] <= 32'b010010_11110_01101_1111111111111111; 	// sw
disk[161] <= 32'b010010_11110_11111_1111111111111101; 	// sw
disk[162] <= 32'b010111_00000000000000000001001110; 	// jal
disk[163] <= 32'b000010_11110_11110_0000000000001001; 	// subi
disk[164] <= 32'b001111_11110_01010_1111111111111001; 	// lw
disk[165] <= 32'b001111_11110_01100_1111111111111001; 	// lw
disk[166] <= 32'b001111_11110_01101_1111111111111111; 	// lw
disk[167] <= 32'b001111_11110_11111_1111111111111101; 	// lw
disk[168] <= 32'b001110_00001_01110_0000000000000000; 	// mov
disk[169] <= 32'b001111_11110_01111_0000000000000000; 	// lw
disk[170] <= 32'b001110_01111_00110_0000000000000000; 	// mov
disk[171] <= 32'b010000_00000_00111_0000000000000011; 	// li
disk[172] <= 32'b010010_11110_01010_1111111111111001; 	// sw
disk[173] <= 32'b010010_11110_01100_1111111111111001; 	// sw
disk[174] <= 32'b010010_11110_01101_1111111111111111; 	// sw
disk[175] <= 32'b010010_11110_01110_1111111111111001; 	// sw
disk[176] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[177] <= 32'b010010_11110_11111_1111111111111101; 	// sw
disk[178] <= 32'b010111_00000000000000000001001110; 	// jal
disk[179] <= 32'b000010_11110_11110_0000000000001001; 	// subi
disk[180] <= 32'b001111_11110_01010_1111111111111001; 	// lw
disk[181] <= 32'b001111_11110_01100_1111111111111001; 	// lw
disk[182] <= 32'b001111_11110_01101_1111111111111111; 	// lw
disk[183] <= 32'b001111_11110_01110_1111111111111001; 	// lw
disk[184] <= 32'b001111_11110_01111_0000000000000000; 	// lw
disk[185] <= 32'b001111_11110_11111_1111111111111101; 	// lw
disk[186] <= 32'b001110_00001_10000_0000000000000000; 	// mov
disk[187] <= 32'b010000_00000_00110_0000000000000001; 	// li
disk[188] <= 32'b100100_00110_00000_0000000000000000; 	// mmuSelect
disk[189] <= 32'b100110_00000000000000000000000000; 	// exec
disk[190] <= 32'b010000_00000_00110_0000000000000010; 	// li
disk[191] <= 32'b100100_00110_00000_0000000000000000; 	// mmuSelect
disk[192] <= 32'b100110_00000000000000000000000000; 	// exec
disk[193] <= 32'b010000_00000_00110_0000000000000011; 	// li
disk[194] <= 32'b100100_00110_00000_0000000000000000; 	// mmuSelect
disk[195] <= 32'b100110_00000000000000000000000000; 	// exec
disk[196] <= 32'b011000_00000000000000000000000000; 	// halt
		
		// PROGRAMA 1
		disk[250] <= 32'b010110_00000000000000000000100001;		// Jump to Main
		disk[251] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[252] <= 32'b010010_11110_00110_1111111111111100; 	// sw
		disk[253] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[254] <= 32'b010010_11110_10100_1111111111111111; 	// sw
		disk[255] <= 32'b010000_00000_10101_0000000000000001; 	// li
		disk[256] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[257] <= 32'b010000_00000_10110_0000000000000000; 	// li
		disk[258] <= 32'b010010_11110_10110_1111111111111101; 	// sw
		disk[259] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[260] <= 32'b001111_11110_01011_1111111111111100; 	// lw
		disk[261] <= 32'b000000_01010_01011_10111_00000_001111; 	// let
		disk[262] <= 32'b010101_10111_00000_0000000000011111; 	// jf
		disk[263] <= 32'b010000_00000_11001_0000000000000001; 	// li
		disk[264] <= 32'b000000_01010_11001_11000_00000_001111; 	// let
		disk[265] <= 32'b010101_11000_00000_0000000000010010; 	// jf
		disk[266] <= 32'b010010_11110_01010_1111111111111110; 	// sw
		disk[267] <= 32'b010110_00000000000000000000011011; 	// j
		disk[268] <= 32'b001111_11110_01100_1111111111111111; 	// lw
		disk[269] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[270] <= 32'b000000_01100_01101_11010_00000_000000; 	// add
		disk[271] <= 32'b010010_11110_11010_1111111111111110; 	// sw
		disk[272] <= 32'b010010_11110_01101_1111111111111111; 	// sw
		disk[273] <= 32'b001111_11110_01100_1111111111111111; 	// lw
		disk[274] <= 32'b001111_11110_01110_1111111111111110; 	// lw
		disk[275] <= 32'b010010_11110_01110_0000000000000000; 	// sw
		disk[276] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[277] <= 32'b000001_01010_11011_0000000000000001; 	// addi
		disk[278] <= 32'b010010_11110_11011_1111111111111101; 	// sw
		disk[279] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[280] <= 32'b010110_00000000000000000000001001; 	// j
		disk[281] <= 32'b001110_01110_00001_0000000000000000; 	// mov
		disk[282] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[283] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[284] <= 32'b010000_00000_10100_0000000000001011; 	// li
		disk[285] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[286] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[287] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[288] <= 32'b010010_11110_01010_0000000000000000; 	// sw
		disk[289] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[290] <= 32'b010111_00000000000000000000000001; 	// jal
		disk[291] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[292] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[293] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[294] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[295] <= 32'b001110_01011_00110_0000000000000000; 	// mov
		disk[296] <= 32'b010000_00000_00111_0000000000000000; 	// li
		disk[297] <= 32'b010100_00000_00110_0000000000000000; 	// out
		disk[298] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[299] <= 32'b100101_11111_00000_0000000000000000; 	// syscall

		// PROGRAMA 2
		disk[300] <= 32'b010110_00000000000000000000011111;		// Jump to Main
		disk[301] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[302] <= 32'b010010_11110_00110_1111111111111100; 	// sw
		disk[303] <= 32'b010010_11110_00111_1111111111111101; 	// sw
		disk[304] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[305] <= 32'b010010_11110_10100_1111111111111110; 	// sw
		disk[306] <= 32'b010000_00000_10101_0000000000000000; 	// li
		disk[307] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[308] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[309] <= 32'b001111_11110_01011_1111111111111101; 	// lw
		disk[310] <= 32'b000000_01010_01011_10110_00000_001110; 	// lt
		disk[311] <= 32'b010101_10110_00000_0000000000011011; 	// jf
		disk[312] <= 32'b001111_11110_01100_1111111111111100; 	// lw
		disk[313] <= 32'b000000_01100_01010_10111_00000_000000; 	// add
		disk[314] <= 32'b001111_10111_10111_0000000000000000; 	// lw
		disk[315] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[316] <= 32'b000000_01101_10111_11000_00000_001110; 	// lt
		disk[317] <= 32'b010101_11000_00000_0000000000010111; 	// jf
		disk[318] <= 32'b000000_01100_01010_11001_00000_000000; 	// add
		disk[319] <= 32'b001111_11001_11001_0000000000000000; 	// lw
		disk[320] <= 32'b010010_11110_11001_0000000000000000; 	// sw
		disk[321] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[322] <= 32'b010010_11110_01010_1111111111111111; 	// sw
		disk[323] <= 32'b000001_01010_11010_0000000000000001; 	// addi
		disk[324] <= 32'b010010_11110_11010_1111111111111110; 	// sw
		disk[325] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[326] <= 32'b010110_00000000000000000000001000; 	// j
		disk[327] <= 32'b001110_01101_00110_0000000000000000; 	// mov
		disk[328] <= 32'b010000_00000_00111_0000000000000001; 	// li
		disk[329] <= 32'b010100_00000_00110_0000000000000001; 	// out
		disk[330] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[331] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[332] <= 32'b010001_11110_01010_1111111111111011; 	// la
		disk[333] <= 32'b010000_00000_10100_0000000000001100; 	// li
		disk[334] <= 32'b010010_01010_10100_0000000000000000; 	// sw
		disk[335] <= 32'b010000_00000_10101_0000000000101001; 	// li
		disk[336] <= 32'b010010_01010_10101_0000000000000001; 	// sw
		disk[337] <= 32'b010000_00000_10110_0000000000010111; 	// li
		disk[338] <= 32'b010010_01010_10110_0000000000000010; 	// sw
		disk[339] <= 32'b010000_00000_10111_0000000001100010; 	// li
		disk[340] <= 32'b010010_01010_10111_0000000000000011; 	// sw
		disk[341] <= 32'b010000_00000_11000_0000000000100001; 	// li
		disk[342] <= 32'b010010_01010_11000_0000000000000100; 	// sw
		disk[343] <= 32'b010000_00000_11001_0000000000010101; 	// li
		disk[344] <= 32'b010010_01010_11001_0000000000000101; 	// sw
		disk[345] <= 32'b010001_11110_00110_1111111111111011; 	// la
		disk[346] <= 32'b010000_00000_00111_0000000000000110; 	// li
		disk[347] <= 32'b010010_11110_11111_1111111111111010; 	// sw
		disk[348] <= 32'b010111_00000000000000000000000001; 	// jal
		disk[349] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[350] <= 32'b001111_11110_11111_1111111111111010; 	// lw
		disk[351] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[352] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[353] <= 32'b100101_11111_00000_0000000000000000; 	// syscall
		
		// PROGRAMA 3
		disk[354] <= 32'b010110_00000000000000000000010011;		// Jump to Main
		disk[355] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[356] <= 32'b010010_11110_00110_1111111111111111; 	// sw
		disk[357] <= 32'b010000_00000_10100_0000000000000001; 	// li
		disk[358] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[359] <= 32'b001111_11110_01010_1111111111111111; 	// lw
		disk[360] <= 32'b010000_00000_10110_0000000000000000; 	// li
		disk[361] <= 32'b000000_01010_10110_10101_00000_010000; 	// gt
		disk[362] <= 32'b010101_10101_00000_0000000000010001; 	// jf
		disk[363] <= 32'b001111_11110_01011_0000000000000000; 	// lw
		disk[364] <= 32'b000000_01011_01010_10111_00000_000010; 	// mul
		disk[365] <= 32'b010010_11110_10111_0000000000000000; 	// sw
		disk[366] <= 32'b001111_11110_01011_0000000000000000; 	// lw
		disk[367] <= 32'b000010_01010_11000_0000000000000001; 	// subi
		disk[368] <= 32'b010010_11110_11000_1111111111111111; 	// sw
		disk[369] <= 32'b001111_11110_01010_1111111111111111; 	// lw
		disk[370] <= 32'b010110_00000000000000000000000101; 	// j
		disk[371] <= 32'b001110_01011_00001_0000000000000000; 	// mov
		disk[372] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[373] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[374] <= 32'b010000_00000_10100_0000000000000111; 	// li
		disk[375] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[376] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[377] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[378] <= 32'b010010_11110_01010_0000000000000000; 	// sw
		disk[379] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[380] <= 32'b010111_00000000000000000000000001; 	// jal
		disk[381] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[382] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[383] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[384] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[385] <= 32'b001110_01011_00110_0000000000000000; 	// mov
		disk[386] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[387] <= 32'b010100_00000_00110_0000000000000010; 	// out
		disk[388] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[389] <= 32'b100101_11111_00000_0000000000000000; 	// syscall
		
	end
endmodule
