module disco_rigido (clk, we, addr, datain, dataout);
	input clk;										// clock
	input we;										// write enable
	input [31:0] addr;							// disk address
	input [31:0] datain;							// data in (to disk)
	
	output reg [31:0] dataout;					// data out (from disk)
	
	localparam DISK_SIZE = 500;				// Tamanho do disco
	reg [31:0] disk [DISK_SIZE-1:0];			// disk cells
	
	always @ (posedge clk) begin
		if (we) disk[addr] <= datain;			// write disk
	end
	
	always @ (negedge clk) begin
		dataout <= disk[addr];
	end

	initial begin
		// SISTEMA OPERACIONAL
		disk[0] <= 32'b010110_00000000000000000000000001;		// Jump to Main
		disk[1] <= 32'b000001_11110_11110_0000000000001010; 	// addi
		disk[2] <= 32'b010000_00000_00110_0000000000011111; 	// li
		disk[3] <= 32'b010000_00000_00111_0000000000000000; 	// li
		disk[4] <= 32'b010010_00000_00110_0000000000000000; 	// sw
		disk[5] <= 32'b010000_00000_00110_0000000001010101; 	// li
		disk[6] <= 32'b010000_00000_00111_0000000000000001; 	// li
		disk[7] <= 32'b010010_00000_00110_0000000000000001; 	// sw
		disk[8] <= 32'b010000_00000_00110_0000000010001011; 	// li
		disk[9] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[10] <= 32'b010010_00000_00110_0000000000000010; 	// sw
		disk[11] <= 32'b010000_00000_00110_0000000011010010; 	// li
		disk[12] <= 32'b010000_00000_00111_0000000000000011; 	// li
		disk[13] <= 32'b010010_00000_00110_0000000000000011; 	// sw
		disk[14] <= 32'b010000_00000_00110_0000000011111110; 	// li
		disk[15] <= 32'b010000_00000_00111_0000000000000100; 	// li
		disk[16] <= 32'b010010_00000_00110_0000000000000100; 	// sw
		disk[17] <= 32'b010011_00000_10100_0000000000000000; 	// in
		disk[18] <= 32'b001110_10100_00110_0000000000000000; 	// mov
		disk[19] <= 32'b010001_00000_10101_0000000000000000; 	// la
		disk[20] <= 32'b000000_00110_10101_10110_00000_000000; 	// add
		disk[21] <= 32'b001111_10110_10110_0000000000000000; 	// lw
		disk[22] <= 32'b001110_10110_10111_0000000000000000; 	// mov
		disk[23] <= 32'b010010_11110_10111_0000000000000000; 	// sw
		disk[24] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[25] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[26] <= 32'b010000_00000_00111_0000000000000000; 	// li
		disk[27] <= 32'b010100_00000_00110_0000000000000000; 	// out
		disk[28] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[29] <= 32'b000000_00110_00000_00000_00000_010010; 	// jr
		disk[30] <= 32'b011000_00000000000000000000000000; 	// halt
		
		// MAIOR ELEMENTO
		disk[31] <= 32'b010110_00000000000000000001000001;		// Jump to Main
		disk[32] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[33] <= 32'b010010_11110_00110_1111111111111100; 	// sw
		disk[34] <= 32'b010010_11110_00111_1111111111111101; 	// sw
		disk[35] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[36] <= 32'b010010_11110_10100_1111111111111110; 	// sw
		disk[37] <= 32'b010000_00000_10101_0000000000000000; 	// li
		disk[38] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[39] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[40] <= 32'b001111_11110_01011_1111111111111101; 	// lw
		disk[41] <= 32'b000000_01010_01011_10110_00000_001110; 	// lt
		disk[42] <= 32'b010101_10110_00000_0000000000111000; 	// jf
		disk[43] <= 32'b001111_11110_01100_1111111111111100; 	// lw
		disk[44] <= 32'b000000_01100_01010_10111_00000_000000; 	// add
		disk[45] <= 32'b001111_10111_10111_0000000000000000; 	// lw
		disk[46] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[47] <= 32'b000000_01101_10111_11000_00000_001110; 	// lt
		disk[48] <= 32'b010101_11000_00000_0000000000110101; 	// jf
		disk[49] <= 32'b000000_01100_01010_11001_00000_000000; 	// add
		disk[50] <= 32'b001111_11001_11001_0000000000000000; 	// lw
		disk[51] <= 32'b010010_11110_11001_0000000000000000; 	// sw
		disk[52] <= 32'b010010_11110_01010_1111111111111111; 	// sw
		disk[53] <= 32'b000001_01010_11010_0000000000000001; 	// addi
		disk[54] <= 32'b010010_11110_11010_1111111111111110; 	// sw
		disk[55] <= 32'b010110_00000000000000000000100111; 	// j
		disk[56] <= 32'b001111_11110_01110_1111111111111111; 	// lw
		disk[57] <= 32'b001110_01110_00110_0000000000000000; 	// mov
		disk[58] <= 32'b010000_00000_00111_0000000000000001; 	// li
		disk[59] <= 32'b010100_00000_00110_0000000000000001; 	// out
		disk[60] <= 32'b001111_11110_01111_0000000000000000; 	// lw
		disk[61] <= 32'b001110_01111_00110_0000000000000000; 	// mov
		disk[62] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[63] <= 32'b010100_00000_00110_0000000000000010; 	// out
		disk[64] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[65] <= 32'b000001_11110_11110_0000000000000110; 	// addi
		disk[66] <= 32'b010001_11110_01010_1111111111111011; 	// la
		disk[67] <= 32'b010000_00000_10100_0000000000001100; 	// li
		disk[68] <= 32'b010010_01010_10100_0000000000000000; 	// sw
		disk[69] <= 32'b010000_00000_10101_0000000000101001; 	// li
		disk[70] <= 32'b010010_01010_10101_0000000000000001; 	// sw
		disk[71] <= 32'b010000_00000_10110_0000000000010111; 	// li
		disk[72] <= 32'b010010_01010_10110_0000000000000010; 	// sw
		disk[73] <= 32'b010000_00000_10111_0000000001100010; 	// li
		disk[74] <= 32'b010010_01010_10111_0000000000000011; 	// sw
		disk[75] <= 32'b010000_00000_11000_0000000000100001; 	// li
		disk[76] <= 32'b010010_01010_11000_0000000000000100; 	// sw
		disk[77] <= 32'b010000_00000_11001_0000000000010101; 	// li
		disk[78] <= 32'b010010_01010_11001_0000000000000101; 	// sw
		disk[79] <= 32'b010001_11110_00110_1111111111111011; 	// la
		disk[80] <= 32'b010000_00000_00111_0000000000000110; 	// li
		disk[81] <= 32'b010111_00000000000000000000100000; 	// jal
		disk[82] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[83] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[84] <= 32'b011000_00000000000000000000000000; 	// halt
		
		// MENOR ELEMENTO
		disk[85] <= 32'b010110_00000000000000000001110111;		// Jump to Main
		disk[86] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[87] <= 32'b010010_11110_00110_1111111111111100; 	// sw
		disk[88] <= 32'b010010_11110_00111_1111111111111101; 	// sw
		disk[89] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[90] <= 32'b010010_11110_10100_1111111111111110; 	// sw
		disk[91] <= 32'b010000_00000_10101_0000000001100011; 	// li
		disk[92] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[93] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[94] <= 32'b001111_11110_01011_1111111111111101; 	// lw
		disk[95] <= 32'b000000_01010_01011_10110_00000_001110; 	// lt
		disk[96] <= 32'b010101_10110_00000_0000000001101110; 	// jf
		disk[97] <= 32'b001111_11110_01100_1111111111111100; 	// lw
		disk[98] <= 32'b000000_01100_01010_10111_00000_000000; 	// add
		disk[99] <= 32'b001111_10111_10111_0000000000000000; 	// lw
		disk[100] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[101] <= 32'b000000_01101_10111_11000_00000_010000; 	// gt
		disk[102] <= 32'b010101_11000_00000_0000000001101011; 	// jf
		disk[103] <= 32'b000000_01100_01010_11001_00000_000000; 	// add
		disk[104] <= 32'b001111_11001_11001_0000000000000000; 	// lw
		disk[105] <= 32'b010010_11110_11001_0000000000000000; 	// sw
		disk[106] <= 32'b010010_11110_01010_1111111111111111; 	// sw
		disk[107] <= 32'b000001_01010_11010_0000000000000001; 	// addi
		disk[108] <= 32'b010010_11110_11010_1111111111111110; 	// sw
		disk[109] <= 32'b010110_00000000000000000001011101; 	// j
		disk[110] <= 32'b001111_11110_01110_1111111111111111; 	// lw
		disk[111] <= 32'b001110_01110_00110_0000000000000000; 	// mov
		disk[112] <= 32'b010000_00000_00111_0000000000000001; 	// li
		disk[113] <= 32'b010100_00000_00110_0000000000000001; 	// out
		disk[114] <= 32'b001111_11110_01111_0000000000000000; 	// lw
		disk[115] <= 32'b001110_01111_00110_0000000000000000; 	// mov
		disk[116] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[117] <= 32'b010100_00000_00110_0000000000000010; 	// out
		disk[118] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[119] <= 32'b000001_11110_11110_0000000000000110; 	// addi
		disk[120] <= 32'b010001_11110_01010_1111111111111011; 	// la
		disk[121] <= 32'b010000_00000_10100_0000000000001011; 	// li
		disk[122] <= 32'b010010_01010_10100_0000000000000000; 	// sw
		disk[123] <= 32'b010000_00000_10101_0000000000101001; 	// li
		disk[124] <= 32'b010010_01010_10101_0000000000000001; 	// sw
		disk[125] <= 32'b010000_00000_10110_0000000000010111; 	// li
		disk[126] <= 32'b010010_01010_10110_0000000000000010; 	// sw
		disk[127] <= 32'b010000_00000_10111_0000000001100010; 	// li
		disk[128] <= 32'b010010_01010_10111_0000000000000011; 	// sw
		disk[129] <= 32'b010000_00000_11000_0000000000100001; 	// li
		disk[130] <= 32'b010010_01010_11000_0000000000000100; 	// sw
		disk[131] <= 32'b010000_00000_11001_0000000000010101; 	// li
		disk[132] <= 32'b010010_01010_11001_0000000000000101; 	// sw
		disk[133] <= 32'b010001_11110_00110_1111111111111011; 	// la
		disk[134] <= 32'b010000_00000_00111_0000000000000110; 	// li
		disk[135] <= 32'b010111_00000000000000000001010110; 	// jal
		disk[136] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[137] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[138] <= 32'b011000_00000000000000000000000000; 	// halt
		
		// SORT
		disk[139] <= 32'b010110_00000000000000000010111001;		// Jump to Main
		disk[140] <= 32'b000001_11110_11110_0000000000001000; 	// addi
		disk[141] <= 32'b010010_11110_00110_1111111111111011; 	// sw
		disk[142] <= 32'b010010_11110_00111_1111111111111100; 	// sw
		disk[143] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[144] <= 32'b010010_11110_10100_1111111111111101; 	// sw
		disk[145] <= 32'b001111_11110_01010_1111111111111100; 	// lw
		disk[146] <= 32'b000010_01010_10101_0000000000000001; 	// subi
		disk[147] <= 32'b001111_11110_01011_1111111111111101; 	// lw
		disk[148] <= 32'b000000_01011_10101_10110_00000_001110; 	// lt
		disk[149] <= 32'b010101_10110_00000_0000000010111000; 	// jf
		disk[150] <= 32'b010010_11110_01011_1111111111111111; 	// sw
		disk[151] <= 32'b000001_01011_10111_0000000000000001; 	// addi
		disk[152] <= 32'b010010_11110_10111_1111111111111110; 	// sw
		disk[153] <= 32'b001111_11110_01100_1111111111111110; 	// lw
		disk[154] <= 32'b000000_01100_01010_11000_00000_001110; 	// lt
		disk[155] <= 32'b010101_11000_00000_0000000010101000; 	// jf
		disk[156] <= 32'b001111_11110_01101_1111111111111011; 	// lw
		disk[157] <= 32'b000000_01101_01100_11001_00000_000000; 	// add
		disk[158] <= 32'b001111_11001_11001_0000000000000000; 	// lw
		disk[159] <= 32'b001111_11110_01110_1111111111111111; 	// lw
		disk[160] <= 32'b000000_01101_01110_11010_00000_000000; 	// add
		disk[161] <= 32'b001111_11010_11010_0000000000000000; 	// lw
		disk[162] <= 32'b000000_11001_11010_11011_00000_001110; 	// lt
		disk[163] <= 32'b010101_11011_00000_0000000010100101; 	// jf
		disk[164] <= 32'b010010_11110_01100_1111111111111111; 	// sw
		disk[165] <= 32'b000001_01100_11100_0000000000000001; 	// addi
		disk[166] <= 32'b010010_11110_11100_1111111111111110; 	// sw
		disk[167] <= 32'b010110_00000000000000000010011001; 	// j
		disk[168] <= 32'b001111_11110_01111_1111111111111111; 	// lw
		disk[169] <= 32'b000000_01011_01111_11101_00000_001101; 	// ne
		disk[170] <= 32'b010101_11101_00000_0000000010110101; 	// jf
		disk[171] <= 32'b000000_01101_01011_10100_00000_000000; 	// add
		disk[172] <= 32'b001111_10100_10100_0000000000000000; 	// lw
		disk[173] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[174] <= 32'b000000_01101_01111_10101_00000_000000; 	// add
		disk[175] <= 32'b001111_10101_10101_0000000000000000; 	// lw
		disk[176] <= 32'b000000_01101_01011_10110_00000_000000; 	// add
		disk[177] <= 32'b010010_10110_10101_0000000000000000; 	// sw
		disk[178] <= 32'b000000_01101_01111_10111_00000_000000; 	// add
		disk[179] <= 32'b001111_11110_10000_0000000000000000; 	// lw
		disk[180] <= 32'b010010_10111_10000_0000000000000000; 	// sw
		disk[181] <= 32'b000001_01011_11000_0000000000000001; 	// addi
		disk[182] <= 32'b010010_11110_11000_1111111111111101; 	// sw
		disk[183] <= 32'b010110_00000000000000000010010001; 	// j
		disk[184] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[185] <= 32'b000001_11110_11110_0000000000000101; 	// addi
		disk[186] <= 32'b010001_11110_01010_1111111111111100; 	// la
		disk[187] <= 32'b010000_00000_10100_0000000000001001; 	// li
		disk[188] <= 32'b010010_01010_10100_0000000000000000; 	// sw
		disk[189] <= 32'b010000_00000_10101_0000000000000110; 	// li
		disk[190] <= 32'b010010_01010_10101_0000000000000001; 	// sw
		disk[191] <= 32'b010000_00000_10110_0000000000001000; 	// li
		disk[192] <= 32'b010010_01010_10110_0000000000000010; 	// sw
		disk[193] <= 32'b010000_00000_10111_0000000000000111; 	// li
		disk[194] <= 32'b010010_01010_10111_0000000000000011; 	// sw
		disk[195] <= 32'b010001_11110_00110_1111111111111100; 	// la
		disk[196] <= 32'b010000_00000_00111_0000000000000100; 	// li
		disk[197] <= 32'b010111_00000000000000000010001100; 	// jal
		disk[198] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[199] <= 32'b000010_11110_11110_0000000000001000; 	// subi
		disk[200] <= 32'b010011_00000_11000_0000000000000000; 	// in
		disk[201] <= 32'b010010_11110_11000_0000000000000000; 	// sw
		disk[202] <= 32'b010001_11110_01100_1111111111111100; 	// la
		disk[203] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[204] <= 32'b000000_01100_01101_11001_00000_000000; 	// add
		disk[205] <= 32'b001111_11001_11001_0000000000000000; 	// lw
		disk[206] <= 32'b001110_11001_00110_0000000000000000; 	// mov
		disk[207] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[208] <= 32'b010100_00000_00110_0000000000000010; 	// out
		disk[209] <= 32'b011000_00000000000000000000000000; 	// halt
		
		// FIBONACCI
		disk[210] <= 32'b010110_00000000000000000011110000;		// Jump to Main
		disk[211] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[212] <= 32'b010010_11110_00110_1111111111111100; 	// sw
		disk[213] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[214] <= 32'b010010_11110_10100_1111111111111111; 	// sw
		disk[215] <= 32'b010000_00000_10101_0000000000000001; 	// li
		disk[216] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[217] <= 32'b010000_00000_10110_0000000000000000; 	// li
		disk[218] <= 32'b010010_11110_10110_1111111111111101; 	// sw
		disk[219] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[220] <= 32'b001111_11110_01011_1111111111111100; 	// lw
		disk[221] <= 32'b000000_01010_01011_10111_00000_001111; 	// let
		disk[222] <= 32'b010101_10111_00000_0000000011101110; 	// jf
		disk[223] <= 32'b010000_00000_11001_0000000000000001; 	// li
		disk[224] <= 32'b000000_01010_11001_11000_00000_001111; 	// let
		disk[225] <= 32'b010101_11000_00000_0000000011100100; 	// jf
		disk[226] <= 32'b010010_11110_01010_1111111111111110; 	// sw
		disk[227] <= 32'b010110_00000000000000000011101011; 	// j
		disk[228] <= 32'b001111_11110_01100_1111111111111111; 	// lw
		disk[229] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[230] <= 32'b000000_01100_01101_11010_00000_000000; 	// add
		disk[231] <= 32'b010010_11110_11010_1111111111111110; 	// sw
		disk[232] <= 32'b010010_11110_01101_1111111111111111; 	// sw
		disk[233] <= 32'b001111_11110_01110_1111111111111110; 	// lw
		disk[234] <= 32'b010010_11110_01110_0000000000000000; 	// sw
		disk[235] <= 32'b000001_01010_11011_0000000000000001; 	// addi
		disk[236] <= 32'b010010_11110_11011_1111111111111101; 	// sw
		disk[237] <= 32'b010110_00000000000000000011011011; 	// j
		disk[238] <= 32'b001110_01110_00001_0000000000000000; 	// mov
		disk[239] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[240] <= 32'b000001_11110_11110_0000000000000001; 	// addi
		disk[241] <= 32'b010011_00000_10100_0000000000000000; 	// in
		disk[242] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[243] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[244] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[245] <= 32'b010010_11110_01010_0000000000000000; 	// sw
		disk[246] <= 32'b010111_00000000000000000011010011; 	// jal
		disk[247] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[248] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[249] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[250] <= 32'b001110_01011_00110_0000000000000000; 	// mov
		disk[251] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[252] <= 32'b010100_00000_00110_0000000000000010; 	// out
		disk[253] <= 32'b011000_00000000000000000000000000; 	// halt
		
		// FATORIAL
		disk[254] <= 32'b010110_00000000000000000100010000;		// Jump to Main
		disk[255] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[256] <= 32'b010010_11110_00110_1111111111111111; 	// sw
		disk[257] <= 32'b010000_00000_10100_0000000000000001; 	// li
		disk[258] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[259] <= 32'b001111_11110_01010_1111111111111111; 	// lw
		disk[260] <= 32'b010000_00000_10110_0000000000000000; 	// li
		disk[261] <= 32'b000000_01010_10110_10101_00000_010000; 	// gt
		disk[262] <= 32'b010101_10101_00000_0000000100001101; 	// jf
		disk[263] <= 32'b001111_11110_01011_0000000000000000; 	// lw
		disk[264] <= 32'b000000_01011_01010_10111_00000_000010; 	// mul
		disk[265] <= 32'b010010_11110_10111_0000000000000000; 	// sw
		disk[266] <= 32'b000010_01010_11000_0000000000000001; 	// subi
		disk[267] <= 32'b010010_11110_11000_1111111111111111; 	// sw
		disk[268] <= 32'b010110_00000000000000000100000011; 	// j
		disk[269] <= 32'b001111_11110_01100_0000000000000000; 	// lw
		disk[270] <= 32'b001110_01100_00001_0000000000000000; 	// mov
		disk[271] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[272] <= 32'b000001_11110_11110_0000000000000001; 	// addi
		disk[273] <= 32'b010011_00000_10100_0000000000000000; 	// in
		disk[274] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[275] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[276] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[277] <= 32'b010010_11110_01010_0000000000000000; 	// sw
		disk[278] <= 32'b010111_00000000000000000011111111; 	// jal
		disk[279] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[280] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[281] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[282] <= 32'b001110_01011_00110_0000000000000000; 	// mov
		disk[283] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[284] <= 32'b010100_00000_00110_0000000000000010; 	// out
		disk[285] <= 32'b011000_00000000000000000000000000; 	// halt
	end
endmodule
