module disco_rigido (clk, we, addr, datain, dataout);
	input clk;										// clock
	input we;										// write enable
	input [31:0] addr;							// disk address
	input [31:0] datain;							// data in (to disk)
	
	output reg [31:0] dataout;					// data out (from disk)
	
	localparam DISK_SIZE = 4096;				// Tamanho do disco
	reg [31:0] disk [DISK_SIZE-1:0];			// disk cells
	
	always @ (posedge clk) begin
		if (we) disk[addr] <= datain;			// write disk
	end
	
	always @ (negedge clk) begin
		dataout <= disk[addr];
	end

	initial begin
		// SISTEMA OPERACIONAL
		disk[0] <= 32'b111100_00000000000000011000010101;		// Jump to Main
		disk[1] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[2] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[3] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[4] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[5] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[6] <= 32'b010110_00001_10000_0000000000000000; 	// ldk
		disk[7] <= 32'b010010_11110_10000_1111111111111111; 	// sw
		disk[8] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[9] <= 32'b001101_00101_10001_0000000000011010; 	// srli
		disk[10] <= 32'b001111_11101_00110_0000000110101010; 	// lw
		disk[11] <= 32'b000000_10001_00110_10010_00000_001101; 	// ne
		disk[12] <= 32'b010101_10010_00000_0000000000010110; 	// jf
		disk[13] <= 32'b001111_11110_00111_0000000000000000; 	// lw
		disk[14] <= 32'b000001_00111_10011_0000000000000001; 	// addi
		disk[15] <= 32'b010010_11110_10011_0000000000000000; 	// sw
		disk[16] <= 32'b001111_11110_00111_0000000000000000; 	// lw
		disk[17] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[18] <= 32'b010110_00001_10100_0000000000000000; 	// ldk
		disk[19] <= 32'b010010_11110_10100_1111111111111111; 	// sw
		disk[20] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[21] <= 32'b111100_00000000000000000000001000; 	// j
		disk[22] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[23] <= 32'b001110_00101_11000_0000000000000000; 	// mov
		disk[24] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[25] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[26] <= 32'b010010_11110_00001_1111111111111111; 	// sw
		disk[27] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[28] <= 32'b010000_00000_10000_0000000000000000; 	// li
		disk[29] <= 32'b000000_00101_10000_01111_00000_001100; 	// eq
		disk[30] <= 32'b010101_01111_00000_0000000000100010; 	// jf
		disk[31] <= 32'b010000_00000_10001_0000000000000001; 	// li
		disk[32] <= 32'b001110_10001_11000_0000000000000000; 	// mov
		disk[33] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[34] <= 32'b010000_00000_10010_0000000000000001; 	// li
		disk[35] <= 32'b010010_11110_10010_0000000000000000; 	// sw
		disk[36] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[37] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[38] <= 32'b000000_00101_10100_10011_00000_010000; 	// gt
		disk[39] <= 32'b010101_10011_00000_0000000000110000; 	// jf
		disk[40] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[41] <= 32'b000011_00110_10101_0000000000000010; 	// muli
		disk[42] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[43] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[44] <= 32'b000010_00101_10110_0000000000000001; 	// subi
		disk[45] <= 32'b010010_11110_10110_1111111111111111; 	// sw
		disk[46] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[47] <= 32'b111100_00000000000000000000100100; 	// j
		disk[48] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[49] <= 32'b001110_00101_11000_0000000000000000; 	// mov
		disk[50] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[51] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[52] <= 32'b010000_00000_00001_0000000000000000; 	// li
		disk[53] <= 32'b010000_00000_00010_0000000000000000; 	// li
		disk[54] <= 32'b010100_00000_00001_0000000000000000; 	// out
		disk[55] <= 32'b010000_00000_00001_0000000000000000; 	// li
		disk[56] <= 32'b010000_00000_00010_0000000000000001; 	// li
		disk[57] <= 32'b010100_00000_00001_0000000000000001; 	// out
		disk[58] <= 32'b010000_00000_00001_0000000000000000; 	// li
		disk[59] <= 32'b010000_00000_00010_0000000000000010; 	// li
		disk[60] <= 32'b010100_00000_00001_0000000000000010; 	// out
		disk[61] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[62] <= 32'b000001_11110_11110_0000000000000110; 	// addi
		disk[63] <= 32'b010001_11101_00101_0000000001000000; 	// la
		disk[64] <= 32'b001111_11101_00110_0000000001011111; 	// lw
		disk[65] <= 32'b000000_00101_00110_01111_00000_000000; 	// add
		disk[66] <= 32'b001111_01111_01111_0000000000000000; 	// lw
		disk[67] <= 32'b000001_01111_10000_0000000000000001; 	// addi
		disk[68] <= 32'b010010_11110_10000_1111111111111110; 	// sw
		disk[69] <= 32'b001111_11110_00111_1111111111111110; 	// lw
		disk[70] <= 32'b001111_11101_01000_0000000011101011; 	// lw
		disk[71] <= 32'b000000_00111_01000_10001_00000_000010; 	// mul
		disk[72] <= 32'b010010_11110_10001_1111111111111111; 	// sw
		disk[73] <= 32'b001111_11101_01001_0000000011101100; 	// lw
		disk[74] <= 32'b000010_01001_10010_0000000000000001; 	// subi
		disk[75] <= 32'b000000_01000_10010_10011_00000_000010; 	// mul
		disk[76] <= 32'b010010_11110_10011_0000000000000000; 	// sw
		disk[77] <= 32'b001111_11101_00101_0000000011101011; 	// lw
		disk[78] <= 32'b001111_11101_00110_0000000011101100; 	// lw
		disk[79] <= 32'b000000_00101_00110_10100_00000_000010; 	// mul
		disk[80] <= 32'b001111_11110_00111_0000000000000000; 	// lw
		disk[81] <= 32'b000000_00111_10100_10101_00000_001110; 	// lt
		disk[82] <= 32'b010101_10101_00000_0000000001100010; 	// jf
		disk[83] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[84] <= 32'b001110_01000_00001_0000000000000000; 	// mov
		disk[85] <= 32'b001111_00001_10110_0000000000000000; 	// lw
		disk[86] <= 32'b010010_11110_10110_1111111111111101; 	// sw
		disk[87] <= 32'b001111_11110_01001_1111111111111101; 	// lw
		disk[88] <= 32'b001110_01001_00001_0000000000000000; 	// mov
		disk[89] <= 32'b001110_00111_00010_0000000000000000; 	// mov
		disk[90] <= 32'b010010_00010_00001_0000000000000000; 	// sw
		disk[91] <= 32'b000001_01000_10111_0000000000000001; 	// addi
		disk[92] <= 32'b010010_11110_10111_1111111111111111; 	// sw
		disk[93] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[94] <= 32'b000001_00111_01111_0000000000000001; 	// addi
		disk[95] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[96] <= 32'b001111_11110_00111_0000000000000000; 	// lw
		disk[97] <= 32'b111100_00000000000000000001001101; 	// j
		disk[98] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[99] <= 32'b000001_11110_11110_0000000000000110; 	// addi
		disk[100] <= 32'b010010_11110_00001_1111111111111101; 	// sw
		disk[101] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[102] <= 32'b000001_00101_01111_0000000000000001; 	// addi
		disk[103] <= 32'b010010_11110_01111_1111111111111101; 	// sw
		disk[104] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[105] <= 32'b001111_11101_00110_0000000011101100; 	// lw
		disk[106] <= 32'b000010_00110_10000_0000000000000001; 	// subi
		disk[107] <= 32'b001111_11101_00111_0000000011101011; 	// lw
		disk[108] <= 32'b000000_00111_10000_10001_00000_000010; 	// mul
		disk[109] <= 32'b010010_11110_10001_1111111111111111; 	// sw
		disk[110] <= 32'b000000_00101_00111_10010_00000_000010; 	// mul
		disk[111] <= 32'b010010_11110_10010_0000000000000000; 	// sw
		disk[112] <= 32'b001111_11101_00101_0000000011101011; 	// lw
		disk[113] <= 32'b001111_11101_00110_0000000011101100; 	// lw
		disk[114] <= 32'b000000_00101_00110_10011_00000_000010; 	// mul
		disk[115] <= 32'b001111_11110_00111_1111111111111111; 	// lw
		disk[116] <= 32'b000000_00111_10011_10100_00000_001110; 	// lt
		disk[117] <= 32'b010101_10100_00000_0000000010000101; 	// jf
		disk[118] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[119] <= 32'b001111_00001_10101_0000000000000000; 	// lw
		disk[120] <= 32'b010010_11110_10101_1111111111111110; 	// sw
		disk[121] <= 32'b001111_11110_01000_1111111111111110; 	// lw
		disk[122] <= 32'b001110_01000_00001_0000000000000000; 	// mov
		disk[123] <= 32'b001111_11110_01001_0000000000000000; 	// lw
		disk[124] <= 32'b001110_01001_00010_0000000000000000; 	// mov
		disk[125] <= 32'b010010_00010_00001_0000000000000000; 	// sw
		disk[126] <= 32'b000001_00111_10110_0000000000000001; 	// addi
		disk[127] <= 32'b010010_11110_10110_1111111111111111; 	// sw
		disk[128] <= 32'b001111_11110_00111_1111111111111111; 	// lw
		disk[129] <= 32'b000001_01001_10111_0000000000000001; 	// addi
		disk[130] <= 32'b010010_11110_10111_0000000000000000; 	// sw
		disk[131] <= 32'b001111_11110_01001_0000000000000000; 	// lw
		disk[132] <= 32'b111100_00000000000000000001110000; 	// j
		disk[133] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[134] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[135] <= 32'b010010_11110_00001_1111111111111111; 	// sw
		disk[136] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[137] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[138] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[139] <= 32'b001111_11101_00110_0000000011101110; 	// lw
		disk[140] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
		disk[141] <= 32'b010101_10000_00000_0000000010011111; 	// jf
		disk[142] <= 32'b010001_11101_00111_0000000110001010; 	// la
		disk[143] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
		disk[144] <= 32'b001111_10001_10001_0000000000000000; 	// lw
		disk[145] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[146] <= 32'b000000_10001_01000_10010_00000_001100; 	// eq
		disk[147] <= 32'b010101_10010_00000_0000000010011010; 	// jf
		disk[148] <= 32'b010001_11101_01001_0000000101110110; 	// la
		disk[149] <= 32'b000000_01001_00101_10011_00000_000000; 	// add
		disk[150] <= 32'b001111_10011_10011_0000000000000000; 	// lw
		disk[151] <= 32'b000010_10011_10100_0000000000000001; 	// subi
		disk[152] <= 32'b001110_10100_11000_0000000000000000; 	// mov
		disk[153] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[154] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[155] <= 32'b000001_00101_10101_0000000000000001; 	// addi
		disk[156] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[157] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[158] <= 32'b111100_00000000000000000010001010; 	// j
		disk[159] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[160] <= 32'b000001_11110_11110_0000000000000101; 	// addi
		disk[161] <= 32'b010010_11110_00001_1111111111111110; 	// sw
		disk[162] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[163] <= 32'b000010_00101_01111_0000000000000001; 	// subi
		disk[164] <= 32'b010010_11101_01111_0000000001011111; 	// sw
		disk[165] <= 32'b010001_11101_00110_0000000000110110; 	// la
		disk[166] <= 32'b001111_11101_00111_0000000001011111; 	// lw
		disk[167] <= 32'b000000_00110_00111_10000_00000_000000; 	// add
		disk[168] <= 32'b001111_10000_10000_0000000000000000; 	// lw
		disk[169] <= 32'b010010_11110_10000_1111111111111111; 	// sw
		disk[170] <= 32'b010001_11101_01000_0000000001001010; 	// la
		disk[171] <= 32'b000000_01000_00111_10001_00000_000000; 	// add
		disk[172] <= 32'b001111_10001_10001_0000000000000000; 	// lw
		disk[173] <= 32'b010010_11110_10001_0000000000000000; 	// sw
		disk[174] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[175] <= 32'b010000_00000_10011_0000000000000000; 	// li
		disk[176] <= 32'b000000_00101_10011_10010_00000_010000; 	// gt
		disk[177] <= 32'b010101_10010_00000_0000000010111110; 	// jf
		disk[178] <= 32'b010001_11101_00110_0000000001101011; 	// la
		disk[179] <= 32'b001111_11110_00111_1111111111111111; 	// lw
		disk[180] <= 32'b000000_00110_00111_10100_00000_000000; 	// add
		disk[181] <= 32'b010000_00000_10101_0000000000000000; 	// li
		disk[182] <= 32'b010010_10100_10101_0000000000000000; 	// sw
		disk[183] <= 32'b000001_00111_10110_0000000000000001; 	// addi
		disk[184] <= 32'b010010_11110_10110_1111111111111111; 	// sw
		disk[185] <= 32'b001111_11110_00111_1111111111111111; 	// lw
		disk[186] <= 32'b000010_00101_10111_0000000000000001; 	// subi
		disk[187] <= 32'b010010_11110_10111_0000000000000000; 	// sw
		disk[188] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[189] <= 32'b111100_00000000000000000010101110; 	// j
		disk[190] <= 32'b010001_11101_00101_0000000110010100; 	// la
		disk[191] <= 32'b001111_11101_00110_0000000001011111; 	// lw
		disk[192] <= 32'b000000_00101_00110_01111_00000_000000; 	// add
		disk[193] <= 32'b010000_00000_10000_0000000000000000; 	// li
		disk[194] <= 32'b010010_01111_10000_0000000000000000; 	// sw
		disk[195] <= 32'b010001_11101_00111_0000000000000100; 	// la
		disk[196] <= 32'b000000_00111_00110_10001_00000_000000; 	// add
		disk[197] <= 32'b010000_00000_10010_0000000000000000; 	// li
		disk[198] <= 32'b010010_10001_10010_0000000000000000; 	// sw
		disk[199] <= 32'b010001_11101_01000_0000000000001110; 	// la
		disk[200] <= 32'b000000_01000_00110_10011_00000_000000; 	// add
		disk[201] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[202] <= 32'b010010_10011_10100_0000000000000000; 	// sw
		disk[203] <= 32'b010001_11101_01001_0000000000011000; 	// la
		disk[204] <= 32'b000000_01001_00110_10101_00000_000000; 	// add
		disk[205] <= 32'b010000_00000_10110_0000000000000000; 	// li
		disk[206] <= 32'b010010_10101_10110_0000000000000000; 	// sw
		disk[207] <= 32'b010001_11101_01010_0000000000100010; 	// la
		disk[208] <= 32'b000000_01010_00110_10111_00000_000000; 	// add
		disk[209] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[210] <= 32'b010010_10111_01111_0000000000000000; 	// sw
		disk[211] <= 32'b010001_11101_01011_0000000000101100; 	// la
		disk[212] <= 32'b000000_01011_00110_10000_00000_000000; 	// add
		disk[213] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[214] <= 32'b010010_10000_10001_0000000000000000; 	// sw
		disk[215] <= 32'b010001_11101_01100_0000000001000000; 	// la
		disk[216] <= 32'b000000_01100_00110_10010_00000_000000; 	// add
		disk[217] <= 32'b010000_00000_10011_0000000000000000; 	// li
		disk[218] <= 32'b010010_10010_10011_0000000000000000; 	// sw
		disk[219] <= 32'b010001_11101_01101_0000000001001010; 	// la
		disk[220] <= 32'b000000_01101_00110_10100_00000_000000; 	// add
		disk[221] <= 32'b010000_00000_10101_0000000000000000; 	// li
		disk[222] <= 32'b010010_10100_10101_0000000000000000; 	// sw
		disk[223] <= 32'b010001_11101_01110_0000000001010100; 	// la
		disk[224] <= 32'b000000_01110_00110_10110_00000_000000; 	// add
		disk[225] <= 32'b010000_00000_10111_0000000000000000; 	// li
		disk[226] <= 32'b010010_10110_10111_0000000000000000; 	// sw
		disk[227] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[228] <= 32'b010010_11101_01111_0000000001011111; 	// sw
		disk[229] <= 32'b001111_11101_00110_0000000001011111; 	// lw
		disk[230] <= 32'b010000_00000_10000_0000001111100111; 	// li
		disk[231] <= 32'b010010_11101_10000_0000000001011110; 	// sw
		disk[232] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[233] <= 32'b000001_11110_11110_0000000000000101; 	// addi
		disk[234] <= 32'b010010_11110_00001_1111111111111110; 	// sw
		disk[235] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[236] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[237] <= 32'b010010_11110_11111_1111111111111101; 	// sw
		disk[238] <= 32'b111110_00000000000000000010000110; 	// jal
		disk[239] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[240] <= 32'b001111_11110_11111_1111111111111101; 	// lw
		disk[241] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[242] <= 32'b010010_11110_00101_1111111111111110; 	// sw
		disk[243] <= 32'b010001_11101_00110_0000000000000100; 	// la
		disk[244] <= 32'b001111_11110_00111_1111111111111110; 	// lw
		disk[245] <= 32'b000000_00110_00111_01111_00000_000000; 	// add
		disk[246] <= 32'b001111_01111_01111_0000000000000000; 	// lw
		disk[247] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[248] <= 32'b000000_01111_10001_10000_00000_001101; 	// ne
		disk[249] <= 32'b010101_10000_00000_0000000100000001; 	// jf
		disk[250] <= 32'b000001_00111_10010_0000000000000001; 	// addi
		disk[251] <= 32'b001110_10010_00001_0000000000000000; 	// mov
		disk[252] <= 32'b010010_11110_11111_1111111111111101; 	// sw
		disk[253] <= 32'b111110_00000000000000000010100000; 	// jal
		disk[254] <= 32'b000010_11110_11110_0000000000000101; 	// subi
		disk[255] <= 32'b001111_11110_11111_1111111111111101; 	// lw
		disk[256] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[257] <= 32'b010001_11101_00101_0000000110000000; 	// la
		disk[258] <= 32'b001111_11110_00110_1111111111111110; 	// lw
		disk[259] <= 32'b000000_00101_00110_10011_00000_000000; 	// add
		disk[260] <= 32'b001111_10011_10011_0000000000000000; 	// lw
		disk[261] <= 32'b010010_11110_10011_1111111111111111; 	// sw
		disk[262] <= 32'b001111_11110_00111_1111111111111111; 	// lw
		disk[263] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[264] <= 32'b010110_00001_10100_0000000000000000; 	// ldk
		disk[265] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[266] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[267] <= 32'b001101_00101_10101_0000000000011010; 	// srli
		disk[268] <= 32'b001111_11101_00110_0000000110101000; 	// lw
		disk[269] <= 32'b000000_10101_00110_10110_00000_001101; 	// ne
		disk[270] <= 32'b010101_10110_00000_0000000100011011; 	// jf
		disk[271] <= 32'b010000_00000_00001_0000000000000000; 	// li
		disk[272] <= 32'b001111_11110_00111_1111111111111111; 	// lw
		disk[273] <= 32'b001110_00111_00010_0000000000000000; 	// mov
		disk[274] <= 32'b010111_00010_00001_0000000000000000; 	// sdk
		disk[275] <= 32'b000001_00111_10111_0000000000000001; 	// addi
		disk[276] <= 32'b010010_11110_10111_1111111111111111; 	// sw
		disk[277] <= 32'b001111_11110_00111_1111111111111111; 	// lw
		disk[278] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[279] <= 32'b010110_00001_01111_0000000000000000; 	// ldk
		disk[280] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[281] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[282] <= 32'b111100_00000000000000000100001010; 	// j
		disk[283] <= 32'b010000_00000_00001_0000000000000000; 	// li
		disk[284] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[285] <= 32'b001110_00101_00010_0000000000000000; 	// mov
		disk[286] <= 32'b010111_00010_00001_0000000000000000; 	// sdk
		disk[287] <= 32'b010001_11101_00110_0000000101110110; 	// la
		disk[288] <= 32'b001111_11110_00111_1111111111111110; 	// lw
		disk[289] <= 32'b000000_00110_00111_10000_00000_000000; 	// add
		disk[290] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[291] <= 32'b010010_10000_10001_0000000000000000; 	// sw
		disk[292] <= 32'b010001_11101_01000_0000000110001010; 	// la
		disk[293] <= 32'b000000_01000_00111_10010_00000_000000; 	// add
		disk[294] <= 32'b010000_00000_10011_0000000000000000; 	// li
		disk[295] <= 32'b010010_10010_10011_0000000000000000; 	// sw
		disk[296] <= 32'b010001_11101_01001_0000000110000000; 	// la
		disk[297] <= 32'b000000_01001_00111_10100_00000_000000; 	// add
		disk[298] <= 32'b010000_00000_10101_0000000000000000; 	// li
		disk[299] <= 32'b010010_10100_10101_0000000000000000; 	// sw
		disk[300] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[301] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[302] <= 32'b010010_11110_00001_1111111111111111; 	// sw
		disk[303] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[304] <= 32'b000010_00101_01111_0000000000000001; 	// subi
		disk[305] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[306] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[307] <= 32'b001111_11101_00110_0000000110101111; 	// lw
		disk[308] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[309] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[310] <= 32'b010011_00000_10000_0000000000000000; 	// in
		disk[311] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[312] <= 32'b010001_11101_00111_0000000110001010; 	// la
		disk[313] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
		disk[314] <= 32'b001111_11110_01000_0000000000000000; 	// lw
		disk[315] <= 32'b010010_10001_01000_0000000000000000; 	// sw
		disk[316] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[317] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[318] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[319] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[320] <= 32'b010000_00000_10000_0000000000000000; 	// li
		disk[321] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[322] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[323] <= 32'b001111_11101_00110_0000000011101110; 	// lw
		disk[324] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
		disk[325] <= 32'b010101_10001_00000_0000000101011111; 	// jf
		disk[326] <= 32'b010001_11101_00111_0000000101110110; 	// la
		disk[327] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
		disk[328] <= 32'b001111_10010_10010_0000000000000000; 	// lw
		disk[329] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[330] <= 32'b000000_10010_10100_10011_00000_001101; 	// ne
		disk[331] <= 32'b010101_10011_00000_0000000101011010; 	// jf
		disk[332] <= 32'b010001_11101_01000_0000000110001010; 	// la
		disk[333] <= 32'b000000_01000_00101_10101_00000_000000; 	// add
		disk[334] <= 32'b001111_10101_10101_0000000000000000; 	// lw
		disk[335] <= 32'b000010_10101_10110_0000000000000001; 	// subi
		disk[336] <= 32'b001110_10110_00001_0000000000000000; 	// mov
		disk[337] <= 32'b010010_11110_11111_1111111111111110; 	// sw
		disk[338] <= 32'b111110_00000000000000000000011001; 	// jal
		disk[339] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[340] <= 32'b001111_11110_11111_1111111111111110; 	// lw
		disk[341] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[342] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[343] <= 32'b000000_00110_00101_10111_00000_000000; 	// add
		disk[344] <= 32'b010010_11110_10111_0000000000000000; 	// sw
		disk[345] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[346] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[347] <= 32'b000001_00101_01111_0000000000000001; 	// addi
		disk[348] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[349] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[350] <= 32'b111100_00000000000000000101000010; 	// j
		disk[351] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[352] <= 32'b001110_00101_11000_0000000000000000; 	// mov
		disk[353] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[354] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[355] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[356] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[357] <= 32'b010000_00000_10000_0000000000000000; 	// li
		disk[358] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[359] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[360] <= 32'b001111_11101_00110_0000000011101110; 	// lw
		disk[361] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
		disk[362] <= 32'b010101_10001_00000_0000000110000100; 	// jf
		disk[363] <= 32'b010001_11101_00111_0000000110010100; 	// la
		disk[364] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
		disk[365] <= 32'b001111_10010_10010_0000000000000000; 	// lw
		disk[366] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[367] <= 32'b000000_10010_10100_10011_00000_001101; 	// ne
		disk[368] <= 32'b010101_10011_00000_0000000101111111; 	// jf
		disk[369] <= 32'b010001_11101_01000_0000000110001010; 	// la
		disk[370] <= 32'b000000_01000_00101_10101_00000_000000; 	// add
		disk[371] <= 32'b001111_10101_10101_0000000000000000; 	// lw
		disk[372] <= 32'b000010_10101_10110_0000000000000001; 	// subi
		disk[373] <= 32'b001110_10110_00001_0000000000000000; 	// mov
		disk[374] <= 32'b010010_11110_11111_1111111111111110; 	// sw
		disk[375] <= 32'b111110_00000000000000000000011001; 	// jal
		disk[376] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[377] <= 32'b001111_11110_11111_1111111111111110; 	// lw
		disk[378] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[379] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[380] <= 32'b000000_00110_00101_10111_00000_000000; 	// add
		disk[381] <= 32'b010010_11110_10111_0000000000000000; 	// sw
		disk[382] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[383] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[384] <= 32'b000001_00101_01111_0000000000000001; 	// addi
		disk[385] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[386] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[387] <= 32'b111100_00000000000000000101100111; 	// j
		disk[388] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[389] <= 32'b001110_00101_11000_0000000000000000; 	// mov
		disk[390] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[391] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[392] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[393] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[394] <= 32'b010000_00000_10000_0000000000000000; 	// li
		disk[395] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[396] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[397] <= 32'b001111_11101_00110_0000000011101110; 	// lw
		disk[398] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
		disk[399] <= 32'b010101_10001_00000_0000000110101001; 	// jf
		disk[400] <= 32'b010001_11101_00111_0000000000000100; 	// la
		disk[401] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
		disk[402] <= 32'b001111_10010_10010_0000000000000000; 	// lw
		disk[403] <= 32'b001111_11101_01000_0000000000000010; 	// lw
		disk[404] <= 32'b000000_10010_01000_10011_00000_001100; 	// eq
		disk[405] <= 32'b010101_10011_00000_0000000110100100; 	// jf
		disk[406] <= 32'b010001_11101_01001_0000000110001010; 	// la
		disk[407] <= 32'b000000_01001_00101_10100_00000_000000; 	// add
		disk[408] <= 32'b001111_10100_10100_0000000000000000; 	// lw
		disk[409] <= 32'b000010_10100_10101_0000000000000001; 	// subi
		disk[410] <= 32'b001110_10101_00001_0000000000000000; 	// mov
		disk[411] <= 32'b010010_11110_11111_1111111111111110; 	// sw
		disk[412] <= 32'b111110_00000000000000000000011001; 	// jal
		disk[413] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[414] <= 32'b001111_11110_11111_1111111111111110; 	// lw
		disk[415] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[416] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[417] <= 32'b000000_00110_00101_10110_00000_000000; 	// add
		disk[418] <= 32'b010010_11110_10110_0000000000000000; 	// sw
		disk[419] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[420] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[421] <= 32'b000001_00101_10111_0000000000000001; 	// addi
		disk[422] <= 32'b010010_11110_10111_1111111111111111; 	// sw
		disk[423] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[424] <= 32'b111100_00000000000000000110001100; 	// j
		disk[425] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[426] <= 32'b001110_00101_11000_0000000000000000; 	// mov
		disk[427] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[428] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[429] <= 32'b010000_00000_01111_0000000000000010; 	// li
		disk[430] <= 32'b010010_11101_01111_0000000101110100; 	// sw
		disk[431] <= 32'b010000_00000_10000_0000000000000001; 	// li
		disk[432] <= 32'b010010_11101_10000_0000000101110101; 	// sw
		disk[433] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[434] <= 32'b000001_11110_11110_0000000000000011; 	// addi
		disk[435] <= 32'b010000_00000_01111_0000000000000001; 	// li
		disk[436] <= 32'b010010_11101_01111_0000000000000000; 	// sw
		disk[437] <= 32'b010000_00000_10000_0000000000000010; 	// li
		disk[438] <= 32'b010010_11101_10000_0000000000000001; 	// sw
		disk[439] <= 32'b010000_00000_10001_0000000000000011; 	// li
		disk[440] <= 32'b010010_11101_10001_0000000000000010; 	// sw
		disk[441] <= 32'b010000_00000_10010_0000000110010100; 	// li
		disk[442] <= 32'b010010_11101_10010_0000000000000011; 	// sw
		disk[443] <= 32'b010000_00000_10011_0000000000000000; 	// li
		disk[444] <= 32'b010010_11110_10011_0000000000000000; 	// sw
		disk[445] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[446] <= 32'b010000_00000_10101_0000000000001010; 	// li
		disk[447] <= 32'b000000_00101_10101_10100_00000_001110; 	// lt
		disk[448] <= 32'b010101_10100_00000_0000000111101001; 	// jf
		disk[449] <= 32'b010001_11101_00110_0000000000000100; 	// la
		disk[450] <= 32'b000000_00110_00101_10110_00000_000000; 	// add
		disk[451] <= 32'b010000_00000_10111_0000000000000000; 	// li
		disk[452] <= 32'b010010_10110_10111_0000000000000000; 	// sw
		disk[453] <= 32'b010001_11101_00111_0000000000001110; 	// la
		disk[454] <= 32'b000000_00111_00101_01111_00000_000000; 	// add
		disk[455] <= 32'b010000_00000_10000_0000000000000000; 	// li
		disk[456] <= 32'b010010_01111_10000_0000000000000000; 	// sw
		disk[457] <= 32'b010001_11101_01000_0000000000011000; 	// la
		disk[458] <= 32'b000000_01000_00101_10001_00000_000000; 	// add
		disk[459] <= 32'b010000_00000_10010_0000000000000000; 	// li
		disk[460] <= 32'b010010_10001_10010_0000000000000000; 	// sw
		disk[461] <= 32'b010001_11101_01001_0000000000100010; 	// la
		disk[462] <= 32'b000000_01001_00101_10011_00000_000000; 	// add
		disk[463] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[464] <= 32'b010010_10011_10100_0000000000000000; 	// sw
		disk[465] <= 32'b010001_11101_01010_0000000000101100; 	// la
		disk[466] <= 32'b000000_01010_00101_10101_00000_000000; 	// add
		disk[467] <= 32'b010000_00000_10110_0000000000000000; 	// li
		disk[468] <= 32'b010010_10101_10110_0000000000000000; 	// sw
		disk[469] <= 32'b010001_11101_01011_0000000001000000; 	// la
		disk[470] <= 32'b000000_01011_00101_10111_00000_000000; 	// add
		disk[471] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[472] <= 32'b010010_10111_01111_0000000000000000; 	// sw
		disk[473] <= 32'b010001_11101_01100_0000000001001010; 	// la
		disk[474] <= 32'b000000_01100_00101_10000_00000_000000; 	// add
		disk[475] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[476] <= 32'b010010_10000_10001_0000000000000000; 	// sw
		disk[477] <= 32'b010001_11101_01101_0000000001010100; 	// la
		disk[478] <= 32'b000000_01101_00101_10010_00000_000000; 	// add
		disk[479] <= 32'b010000_00000_10011_0000000000000000; 	// li
		disk[480] <= 32'b010010_10010_10011_0000000000000000; 	// sw
		disk[481] <= 32'b010001_11101_01110_0000000001100000; 	// la
		disk[482] <= 32'b000000_01110_00101_10100_00000_000000; 	// add
		disk[483] <= 32'b010000_00000_10101_0000000000000000; 	// li
		disk[484] <= 32'b010010_10100_10101_0000000000000000; 	// sw
		disk[485] <= 32'b000001_00101_10110_0000000000000001; 	// addi
		disk[486] <= 32'b010010_11110_10110_0000000000000000; 	// sw
		disk[487] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[488] <= 32'b111100_00000000000000000110111101; 	// j
		disk[489] <= 32'b010000_00000_10111_0000000000000000; 	// li
		disk[490] <= 32'b010010_11101_10111_0000000001101010; 	// sw
		disk[491] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[492] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[493] <= 32'b010000_00000_01111_0000000000100000; 	// li
		disk[494] <= 32'b010010_11101_01111_0000000011101011; 	// sw
		disk[495] <= 32'b010000_00000_10000_0000000010000000; 	// li
		disk[496] <= 32'b010010_11101_10000_0000000011101100; 	// sw
		disk[497] <= 32'b010000_00000_10001_0000000001100100; 	// li
		disk[498] <= 32'b010010_11101_10001_0000000011101101; 	// sw
		disk[499] <= 32'b010000_00000_10010_0000000000001010; 	// li
		disk[500] <= 32'b010010_11101_10010_0000000011101110; 	// sw
		disk[501] <= 32'b010000_00000_10011_0000001111100111; 	// li
		disk[502] <= 32'b010010_11101_10011_0000000001011110; 	// sw
		disk[503] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[504] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[505] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[506] <= 32'b010010_11101_01111_0000000110101011; 	// sw
		disk[507] <= 32'b010000_00000_10000_0000000000000001; 	// li
		disk[508] <= 32'b010010_11101_10000_0000000110101100; 	// sw
		disk[509] <= 32'b010000_00000_10001_0000000000000010; 	// li
		disk[510] <= 32'b010010_11101_10001_0000000110101101; 	// sw
		disk[511] <= 32'b010000_00000_10010_0000000000000011; 	// li
		disk[512] <= 32'b010010_11101_10010_0000000110101110; 	// sw
		disk[513] <= 32'b010000_00000_10011_0000000000000100; 	// li
		disk[514] <= 32'b010010_11101_10011_0000000110101111; 	// sw
		disk[515] <= 32'b010000_00000_10100_0000000000000101; 	// li
		disk[516] <= 32'b010010_11101_10100_0000000110110000; 	// sw
		disk[517] <= 32'b010000_00000_10101_0000000000000110; 	// li
		disk[518] <= 32'b010010_11101_10101_0000000110110001; 	// sw
		disk[519] <= 32'b010000_00000_10110_0000000000000111; 	// li
		disk[520] <= 32'b010010_11101_10110_0000000110110010; 	// sw
		disk[521] <= 32'b010000_00000_10111_0000000000001000; 	// li
		disk[522] <= 32'b010010_11101_10111_0000000110110011; 	// sw
		disk[523] <= 32'b010000_00000_01111_0000000000001001; 	// li
		disk[524] <= 32'b010010_11101_01111_0000000110110100; 	// sw
		disk[525] <= 32'b010000_00000_10000_0000000000001010; 	// li
		disk[526] <= 32'b010010_11101_10000_0000000110110101; 	// sw
		disk[527] <= 32'b010000_00000_10001_0000000000001011; 	// li
		disk[528] <= 32'b010010_11101_10001_0000000110110110; 	// sw
		disk[529] <= 32'b010000_00000_10010_0000000000001100; 	// li
		disk[530] <= 32'b010010_11101_10010_0000000110110111; 	// sw
		disk[531] <= 32'b010000_00000_10011_0000000000001101; 	// li
		disk[532] <= 32'b010010_11101_10011_0000000110111000; 	// sw
		disk[533] <= 32'b010000_00000_10100_0000000000001110; 	// li
		disk[534] <= 32'b010010_11101_10100_0000000110111001; 	// sw
		disk[535] <= 32'b010000_00000_10101_0000000000001111; 	// li
		disk[536] <= 32'b010010_11101_10101_0000000110111010; 	// sw
		disk[537] <= 32'b010000_00000_10110_0000000000010000; 	// li
		disk[538] <= 32'b010010_11101_10110_0000000110111011; 	// sw
		disk[539] <= 32'b010000_00000_10111_0000000000011110; 	// li
		disk[540] <= 32'b010010_11101_10111_0000000110111100; 	// sw
		disk[541] <= 32'b001111_11101_00101_0000000110101011; 	// lw
		disk[542] <= 32'b010010_11101_00101_0000000110111101; 	// sw
		disk[543] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[544] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[545] <= 32'b010000_00000_01111_0000111111111111; 	// li
		disk[546] <= 32'b010010_11101_01111_0000000011110000; 	// sw
		disk[547] <= 32'b010000_00000_10000_0000000000011111; 	// li
		disk[548] <= 32'b010010_11101_10000_0000000110101000; 	// sw
		disk[549] <= 32'b010000_00000_10001_0000000000111101; 	// li
		disk[550] <= 32'b010010_11101_10001_0000000110101001; 	// sw
		disk[551] <= 32'b010000_00000_10010_0000000000111111; 	// li
		disk[552] <= 32'b010010_11101_10010_0000000110101010; 	// sw
		disk[553] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[554] <= 32'b000001_11110_11110_0000000000000101; 	// addi
		disk[555] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[556] <= 32'b010010_11110_01111_1111111111111110; 	// sw
		disk[557] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[558] <= 32'b001111_11101_00110_0000000011101100; 	// lw
		disk[559] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
		disk[560] <= 32'b010101_10000_00000_0000001000111101; 	// jf
		disk[561] <= 32'b010001_11101_00111_0000000001101011; 	// la
		disk[562] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
		disk[563] <= 32'b010000_00000_10010_0000000000000000; 	// li
		disk[564] <= 32'b010010_10001_10010_0000000000000000; 	// sw
		disk[565] <= 32'b010001_11101_01000_0000000011110100; 	// la
		disk[566] <= 32'b000000_01000_00101_10011_00000_000000; 	// add
		disk[567] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[568] <= 32'b010010_10011_10100_0000000000000000; 	// sw
		disk[569] <= 32'b000001_00101_10101_0000000000000001; 	// addi
		disk[570] <= 32'b010010_11110_10101_1111111111111110; 	// sw
		disk[571] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[572] <= 32'b111100_00000000000000001000101101; 	// j
		disk[573] <= 32'b010010_11110_11111_1111111111111101; 	// sw
		disk[574] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[575] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[576] <= 32'b001111_11110_11111_1111111111111101; 	// lw
		disk[577] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[578] <= 32'b010010_11110_00101_0000000000000000; 	// sw
		disk[579] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[580] <= 32'b000001_00110_10110_0000000000000001; 	// addi
		disk[581] <= 32'b010010_11101_10110_0000000011101111; 	// sw
		disk[582] <= 32'b001111_11101_00111_0000000011101011; 	// lw
		disk[583] <= 32'b000000_00110_00111_10111_00000_000011; 	// div
		disk[584] <= 32'b010010_11110_10111_1111111111111111; 	// sw
		disk[585] <= 32'b000000_00110_00111_01111_00000_000100; 	// mod
		disk[586] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[587] <= 32'b000000_01111_10001_10000_00000_010000; 	// gt
		disk[588] <= 32'b010101_10000_00000_0000001001010001; 	// jf
		disk[589] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[590] <= 32'b000001_01000_10010_0000000000000001; 	// addi
		disk[591] <= 32'b010010_11110_10010_1111111111111111; 	// sw
		disk[592] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[593] <= 32'b010000_00000_10011_0000000000000000; 	// li
		disk[594] <= 32'b010010_11110_10011_1111111111111110; 	// sw
		disk[595] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[596] <= 32'b001111_11110_00110_1111111111111111; 	// lw
		disk[597] <= 32'b000000_00101_00110_10100_00000_001110; 	// lt
		disk[598] <= 32'b010101_10100_00000_0000001001011111; 	// jf
		disk[599] <= 32'b010001_11101_00111_0000000001101011; 	// la
		disk[600] <= 32'b000000_00111_00101_10101_00000_000000; 	// add
		disk[601] <= 32'b010000_00000_10110_0000000000000001; 	// li
		disk[602] <= 32'b010010_10101_10110_0000000000000000; 	// sw
		disk[603] <= 32'b000001_00101_10111_0000000000000001; 	// addi
		disk[604] <= 32'b010010_11110_10111_1111111111111110; 	// sw
		disk[605] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[606] <= 32'b111100_00000000000000001001010011; 	// j
		disk[607] <= 32'b001110_11110_01111_0000000000000000; 	// mov
		disk[608] <= 32'b001111_11101_00101_0000000011101011; 	// lw
		disk[609] <= 32'b000000_01111_00101_10000_00000_000011; 	// div
		disk[610] <= 32'b010010_11110_10000_1111111111111111; 	// sw
		disk[611] <= 32'b001110_11110_10001_0000000000000000; 	// mov
		disk[612] <= 32'b000000_10001_00101_10010_00000_000100; 	// mod
		disk[613] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[614] <= 32'b000000_10010_10100_10011_00000_010000; 	// gt
		disk[615] <= 32'b010101_10011_00000_0000001001101100; 	// jf
		disk[616] <= 32'b001111_11110_00110_1111111111111111; 	// lw
		disk[617] <= 32'b000001_00110_10101_0000000000000001; 	// addi
		disk[618] <= 32'b010010_11110_10101_1111111111111111; 	// sw
		disk[619] <= 32'b001111_11110_00110_1111111111111111; 	// lw
		disk[620] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[621] <= 32'b000001_00101_10110_0000000000000001; 	// addi
		disk[622] <= 32'b010010_11110_10110_1111111111111111; 	// sw
		disk[623] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[624] <= 32'b010000_00000_10111_0000000000000000; 	// li
		disk[625] <= 32'b010010_11110_10111_1111111111111110; 	// sw
		disk[626] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[627] <= 32'b001111_11110_00110_1111111111111111; 	// lw
		disk[628] <= 32'b000000_00101_00110_01111_00000_001110; 	// lt
		disk[629] <= 32'b010101_01111_00000_0000001001111110; 	// jf
		disk[630] <= 32'b010001_11101_00111_0000000011110100; 	// la
		disk[631] <= 32'b000000_00111_00101_10000_00000_000000; 	// add
		disk[632] <= 32'b010000_00000_10001_0000000000000001; 	// li
		disk[633] <= 32'b010010_10000_10001_0000000000000000; 	// sw
		disk[634] <= 32'b000001_00101_10010_0000000000000001; 	// addi
		disk[635] <= 32'b010010_11110_10010_1111111111111110; 	// sw
		disk[636] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[637] <= 32'b111100_00000000000000001001110010; 	// j
		disk[638] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[639] <= 32'b001111_11101_00110_0000000011101011; 	// lw
		disk[640] <= 32'b000000_00101_00110_10011_00000_000010; 	// mul
		disk[641] <= 32'b010010_11101_10011_0000000011110001; 	// sw
		disk[642] <= 32'b001111_11101_00111_0000000011101100; 	// lw
		disk[643] <= 32'b000010_00111_10100_0000000000000001; 	// subi
		disk[644] <= 32'b010001_11101_01000_0000000011110100; 	// la
		disk[645] <= 32'b000000_01000_10100_10101_00000_000000; 	// add
		disk[646] <= 32'b010000_00000_10110_0000000000000001; 	// li
		disk[647] <= 32'b010010_10101_10110_0000000000000000; 	// sw
		disk[648] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[649] <= 32'b000001_11110_11110_0000000000000101; 	// addi
		disk[650] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[651] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[652] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[653] <= 32'b001111_11101_00110_0000000011101110; 	// lw
		disk[654] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
		disk[655] <= 32'b010101_10000_00000_0000001010101000; 	// jf
		disk[656] <= 32'b010001_11101_00111_0000000101110110; 	// la
		disk[657] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
		disk[658] <= 32'b010000_00000_10010_0000000000000000; 	// li
		disk[659] <= 32'b010010_10001_10010_0000000000000000; 	// sw
		disk[660] <= 32'b010001_11101_01000_0000000110000000; 	// la
		disk[661] <= 32'b000000_01000_00101_10011_00000_000000; 	// add
		disk[662] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[663] <= 32'b010010_10011_10100_0000000000000000; 	// sw
		disk[664] <= 32'b010001_11101_01001_0000000110001010; 	// la
		disk[665] <= 32'b000000_01001_00101_10101_00000_000000; 	// add
		disk[666] <= 32'b010000_00000_10110_0000000000000000; 	// li
		disk[667] <= 32'b010010_10101_10110_0000000000000000; 	// sw
		disk[668] <= 32'b010001_11101_01010_0000000110010100; 	// la
		disk[669] <= 32'b000000_01010_00101_10111_00000_000000; 	// add
		disk[670] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[671] <= 32'b010010_10111_01111_0000000000000000; 	// sw
		disk[672] <= 32'b010001_11101_01011_0000000110011110; 	// la
		disk[673] <= 32'b000000_01011_00101_10000_00000_000000; 	// add
		disk[674] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[675] <= 32'b010010_10000_10001_0000000000000000; 	// sw
		disk[676] <= 32'b000001_00101_10010_0000000000000001; 	// addi
		disk[677] <= 32'b010010_11110_10010_1111111111111111; 	// sw
		disk[678] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[679] <= 32'b111100_00000000000000001010001100; 	// j
		disk[680] <= 32'b001111_11101_00101_0000000011101111; 	// lw
		disk[681] <= 32'b010010_11110_00101_1111111111111110; 	// sw
		disk[682] <= 32'b010000_00000_10011_0000000000000000; 	// li
		disk[683] <= 32'b010010_11110_10011_1111111111111111; 	// sw
		disk[684] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[685] <= 32'b001111_11101_00110_0000000011110000; 	// lw
		disk[686] <= 32'b000000_00101_00110_10100_00000_001110; 	// lt
		disk[687] <= 32'b010101_10100_00000_0000001011001101; 	// jf
		disk[688] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[689] <= 32'b010110_00001_10101_0000000000000000; 	// ldk
		disk[690] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[691] <= 32'b001111_11110_00111_0000000000000000; 	// lw
		disk[692] <= 32'b001101_00111_10110_0000000000011010; 	// srli
		disk[693] <= 32'b001111_11101_01000_0000000110101001; 	// lw
		disk[694] <= 32'b000000_10110_01000_10111_00000_001100; 	// eq
		disk[695] <= 32'b010101_10111_00000_0000001011001000; 	// jf
		disk[696] <= 32'b001111_11110_01001_1111111111111111; 	// lw
		disk[697] <= 32'b000001_01001_01111_0000000000000001; 	// addi
		disk[698] <= 32'b010001_11101_01010_0000000101110110; 	// la
		disk[699] <= 32'b000000_01010_01001_10000_00000_000000; 	// add
		disk[700] <= 32'b010010_10000_01111_0000000000000000; 	// sw
		disk[701] <= 32'b000000_01010_01001_10001_00000_000000; 	// add
		disk[702] <= 32'b001111_10001_10001_0000000000000000; 	// lw
		disk[703] <= 32'b010001_11101_01011_0000000110001010; 	// la
		disk[704] <= 32'b000000_01011_01001_10010_00000_000000; 	// add
		disk[705] <= 32'b010010_10010_10001_0000000000000000; 	// sw
		disk[706] <= 32'b010001_11101_01100_0000000110000000; 	// la
		disk[707] <= 32'b000000_01100_01001_10011_00000_000000; 	// add
		disk[708] <= 32'b010010_10011_00101_0000000000000000; 	// sw
		disk[709] <= 32'b000001_01001_10100_0000000000000001; 	// addi
		disk[710] <= 32'b010010_11110_10100_1111111111111111; 	// sw
		disk[711] <= 32'b001111_11110_01001_1111111111111111; 	// lw
		disk[712] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[713] <= 32'b000001_00101_10101_0000000000000001; 	// addi
		disk[714] <= 32'b010010_11110_10101_1111111111111110; 	// sw
		disk[715] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[716] <= 32'b111100_00000000000000001010101100; 	// j
		disk[717] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[718] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[719] <= 32'b010010_11110_11111_0000000000000000; 	// sw
		disk[720] <= 32'b111110_00000000000000000110110010; 	// jal
		disk[721] <= 32'b000010_11110_11110_0000000000000011; 	// subi
		disk[722] <= 32'b001111_11110_11111_0000000000000000; 	// lw
		disk[723] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[724] <= 32'b010010_11110_11111_0000000000000000; 	// sw
		disk[725] <= 32'b111110_00000000000000000111101100; 	// jal
		disk[726] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[727] <= 32'b001111_11110_11111_0000000000000000; 	// lw
		disk[728] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[729] <= 32'b010010_11110_11111_0000000000000000; 	// sw
		disk[730] <= 32'b111110_00000000000000000111111000; 	// jal
		disk[731] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[732] <= 32'b001111_11110_11111_0000000000000000; 	// lw
		disk[733] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[734] <= 32'b010010_11110_11111_0000000000000000; 	// sw
		disk[735] <= 32'b111110_00000000000000001000100000; 	// jal
		disk[736] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[737] <= 32'b001111_11110_11111_0000000000000000; 	// lw
		disk[738] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[739] <= 32'b010010_11110_11111_0000000000000000; 	// sw
		disk[740] <= 32'b111110_00000000000000001000101010; 	// jal
		disk[741] <= 32'b000010_11110_11110_0000000000000101; 	// subi
		disk[742] <= 32'b001111_11110_11111_0000000000000000; 	// lw
		disk[743] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[744] <= 32'b010010_11110_11111_0000000000000000; 	// sw
		disk[745] <= 32'b111110_00000000000000001010001001; 	// jal
		disk[746] <= 32'b000010_11110_11110_0000000000000101; 	// subi
		disk[747] <= 32'b001111_11110_11111_0000000000000000; 	// lw
		disk[748] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[749] <= 32'b010010_11110_11111_0000000000000000; 	// sw
		disk[750] <= 32'b111110_00000000000000000110101100; 	// jal
		disk[751] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[752] <= 32'b001111_11110_11111_0000000000000000; 	// lw
		disk[753] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[754] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[755] <= 32'b000001_11110_11110_0000000000000110; 	// addi
		disk[756] <= 32'b010010_11110_00001_1111111111111101; 	// sw
		disk[757] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[758] <= 32'b001111_11101_00110_0000000011101011; 	// lw
		disk[759] <= 32'b000000_00101_00110_01111_00000_000011; 	// div
		disk[760] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[761] <= 32'b000000_00101_00110_10000_00000_000100; 	// mod
		disk[762] <= 32'b010000_00000_10010_0000000000000000; 	// li
		disk[763] <= 32'b000000_10000_10010_10001_00000_010000; 	// gt
		disk[764] <= 32'b010101_10001_00000_0000001100000001; 	// jf
		disk[765] <= 32'b001111_11110_00111_1111111111111111; 	// lw
		disk[766] <= 32'b000001_00111_10011_0000000000000001; 	// addi
		disk[767] <= 32'b010010_11110_10011_1111111111111111; 	// sw
		disk[768] <= 32'b001111_11110_00111_1111111111111111; 	// lw
		disk[769] <= 32'b010001_11101_00101_0000000001001010; 	// la
		disk[770] <= 32'b001111_11101_00110_0000000001011111; 	// lw
		disk[771] <= 32'b000000_00101_00110_10100_00000_000000; 	// add
		disk[772] <= 32'b001111_11110_00111_1111111111111111; 	// lw
		disk[773] <= 32'b010010_10100_00111_0000000000000000; 	// sw
		disk[774] <= 32'b010000_00000_10101_0000000000000000; 	// li
		disk[775] <= 32'b010010_11110_10101_1111111111111110; 	// sw
		disk[776] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[777] <= 32'b001111_11101_00110_0000000011101100; 	// lw
		disk[778] <= 32'b000000_00101_00110_10110_00000_001110; 	// lt
		disk[779] <= 32'b010101_10110_00000_0000001100101011; 	// jf
		disk[780] <= 32'b010001_11101_00111_0000000001101011; 	// la
		disk[781] <= 32'b000000_00111_00101_10111_00000_000000; 	// add
		disk[782] <= 32'b001111_10111_10111_0000000000000000; 	// lw
		disk[783] <= 32'b010000_00000_10000_0000000000000000; 	// li
		disk[784] <= 32'b000000_10111_10000_01111_00000_001100; 	// eq
		disk[785] <= 32'b010101_01111_00000_0000001100100110; 	// jf
		disk[786] <= 32'b010010_11110_00101_0000000000000000; 	// sw
		disk[787] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[788] <= 32'b010000_00000_10010_0000000000000000; 	// li
		disk[789] <= 32'b000000_00101_10010_10001_00000_010000; 	// gt
		disk[790] <= 32'b010101_10001_00000_0000001100100011; 	// jf
		disk[791] <= 32'b010001_11101_00110_0000000001101011; 	// la
		disk[792] <= 32'b001111_11110_00111_1111111111111110; 	// lw
		disk[793] <= 32'b000000_00110_00111_10011_00000_000000; 	// add
		disk[794] <= 32'b010000_00000_10100_0000000000000001; 	// li
		disk[795] <= 32'b010010_10011_10100_0000000000000000; 	// sw
		disk[796] <= 32'b000010_00101_10101_0000000000000001; 	// subi
		disk[797] <= 32'b010010_11110_10101_1111111111111111; 	// sw
		disk[798] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[799] <= 32'b000001_00111_10110_0000000000000001; 	// addi
		disk[800] <= 32'b010010_11110_10110_1111111111111110; 	// sw
		disk[801] <= 32'b001111_11110_00111_1111111111111110; 	// lw
		disk[802] <= 32'b111100_00000000000000001100010011; 	// j
		disk[803] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[804] <= 32'b001110_00101_11000_0000000000000000; 	// mov
		disk[805] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[806] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[807] <= 32'b000001_00101_10111_0000000000000001; 	// addi
		disk[808] <= 32'b010010_11110_10111_1111111111111110; 	// sw
		disk[809] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[810] <= 32'b111100_00000000000000001100001000; 	// j
		disk[811] <= 32'b001111_11101_00101_0000000011101101; 	// lw
		disk[812] <= 32'b001110_00101_11000_0000000000000000; 	// mov
		disk[813] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[814] <= 32'b000001_11110_11110_0000000000000101; 	// addi
		disk[815] <= 32'b010001_11101_00101_0000000000011000; 	// la
		disk[816] <= 32'b001111_11101_00110_0000000001011111; 	// lw
		disk[817] <= 32'b000000_00101_00110_01111_00000_000000; 	// add
		disk[818] <= 32'b001111_01111_01111_0000000000000000; 	// lw
		disk[819] <= 32'b001111_11101_00111_0000000011101011; 	// lw
		disk[820] <= 32'b000000_01111_00111_10000_00000_000011; 	// div
		disk[821] <= 32'b000001_10000_10001_0000000000000001; 	// addi
		disk[822] <= 32'b010010_11110_10001_1111111111111111; 	// sw
		disk[823] <= 32'b000000_00101_00110_10010_00000_000000; 	// add
		disk[824] <= 32'b001111_10010_10010_0000000000000000; 	// lw
		disk[825] <= 32'b000000_10010_00111_10011_00000_000100; 	// mod
		disk[826] <= 32'b010000_00000_10101_0000000000000000; 	// li
		disk[827] <= 32'b000000_10011_10101_10100_00000_010000; 	// gt
		disk[828] <= 32'b010101_10100_00000_0000001101000001; 	// jf
		disk[829] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[830] <= 32'b000001_01000_10110_0000000000000001; 	// addi
		disk[831] <= 32'b010010_11110_10110_1111111111111111; 	// sw
		disk[832] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[833] <= 32'b001111_11101_00101_0000000011101100; 	// lw
		disk[834] <= 32'b000010_00101_10111_0000000000000001; 	// subi
		disk[835] <= 32'b010010_11110_10111_1111111111111110; 	// sw
		disk[836] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[837] <= 32'b010000_00000_10000_0000000000000000; 	// li
		disk[838] <= 32'b000000_00101_10000_01111_00000_010000; 	// gt
		disk[839] <= 32'b010101_01111_00000_0000001101100111; 	// jf
		disk[840] <= 32'b010001_11101_00110_0000000011110100; 	// la
		disk[841] <= 32'b000000_00110_00101_10001_00000_000000; 	// add
		disk[842] <= 32'b001111_10001_10001_0000000000000000; 	// lw
		disk[843] <= 32'b010000_00000_10011_0000000000000000; 	// li
		disk[844] <= 32'b000000_10001_10011_10010_00000_001100; 	// eq
		disk[845] <= 32'b010101_10010_00000_0000001101100010; 	// jf
		disk[846] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[847] <= 32'b010000_00000_10101_0000000000000000; 	// li
		disk[848] <= 32'b000000_00101_10101_10100_00000_010000; 	// gt
		disk[849] <= 32'b010101_10100_00000_0000001101011111; 	// jf
		disk[850] <= 32'b001111_11110_00110_1111111111111110; 	// lw
		disk[851] <= 32'b010010_11110_00110_0000000000000000; 	// sw
		disk[852] <= 32'b010001_11101_00111_0000000011110100; 	// la
		disk[853] <= 32'b000000_00111_00110_10110_00000_000000; 	// add
		disk[854] <= 32'b010000_00000_10111_0000000000000001; 	// li
		disk[855] <= 32'b010010_10110_10111_0000000000000000; 	// sw
		disk[856] <= 32'b000010_00101_01111_0000000000000001; 	// subi
		disk[857] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[858] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[859] <= 32'b000010_00110_10000_0000000000000001; 	// subi
		disk[860] <= 32'b010010_11110_10000_1111111111111110; 	// sw
		disk[861] <= 32'b001111_11110_00110_1111111111111110; 	// lw
		disk[862] <= 32'b111100_00000000000000001101001110; 	// j
		disk[863] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[864] <= 32'b001110_00101_11000_0000000000000000; 	// mov
		disk[865] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[866] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[867] <= 32'b000010_00101_10001_0000000000000001; 	// subi
		disk[868] <= 32'b010010_11110_10001_1111111111111110; 	// sw
		disk[869] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[870] <= 32'b111100_00000000000000001101000100; 	// j
		disk[871] <= 32'b001111_11101_00101_0000000011101101; 	// lw
		disk[872] <= 32'b001110_00101_11000_0000000000000000; 	// mov
		disk[873] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[874] <= 32'b000001_11110_11110_0000000000000011; 	// addi
		disk[875] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[876] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[877] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[878] <= 32'b001111_11101_00110_0000000011101110; 	// lw
		disk[879] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
		disk[880] <= 32'b010101_10000_00000_0000001101111110; 	// jf
		disk[881] <= 32'b010001_11101_00111_0000000000000100; 	// la
		disk[882] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
		disk[883] <= 32'b001111_10001_10001_0000000000000000; 	// lw
		disk[884] <= 32'b001111_11101_01000_0000000000000010; 	// lw
		disk[885] <= 32'b000000_10001_01000_10010_00000_001100; 	// eq
		disk[886] <= 32'b010101_10010_00000_0000001101111001; 	// jf
		disk[887] <= 32'b001110_00101_11000_0000000000000000; 	// mov
		disk[888] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[889] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[890] <= 32'b000001_00101_10011_0000000000000001; 	// addi
		disk[891] <= 32'b010010_11110_10011_0000000000000000; 	// sw
		disk[892] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[893] <= 32'b111100_00000000000000001101101101; 	// j
		disk[894] <= 32'b001111_11101_00101_0000000000000011; 	// lw
		disk[895] <= 32'b001110_00101_11000_0000000000000000; 	// mov
		disk[896] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[897] <= 32'b000001_11110_11110_0000000000000101; 	// addi
		disk[898] <= 32'b010010_11110_00001_1111111111111110; 	// sw
		disk[899] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[900] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[901] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[902] <= 32'b001111_11101_00110_0000000011101110; 	// lw
		disk[903] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
		disk[904] <= 32'b010101_10000_00000_0000001110011001; 	// jf
		disk[905] <= 32'b010001_11101_00111_0000000001100000; 	// la
		disk[906] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
		disk[907] <= 32'b001111_10001_10001_0000000000000000; 	// lw
		disk[908] <= 32'b001111_11110_01000_1111111111111110; 	// lw
		disk[909] <= 32'b000000_10001_01000_10010_00000_001100; 	// eq
		disk[910] <= 32'b010101_10010_00000_0000001110010100; 	// jf
		disk[911] <= 32'b000000_00111_00101_10011_00000_000000; 	// add
		disk[912] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[913] <= 32'b010010_10011_10100_0000000000000000; 	// sw
		disk[914] <= 32'b000001_00101_10101_0000000000000001; 	// addi
		disk[915] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[916] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[917] <= 32'b000001_00101_10110_0000000000000001; 	// addi
		disk[918] <= 32'b010010_11110_10110_1111111111111111; 	// sw
		disk[919] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[920] <= 32'b111100_00000000000000001110000101; 	// j
		disk[921] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[922] <= 32'b001111_11101_00110_0000000011101110; 	// lw
		disk[923] <= 32'b000000_00101_00110_10111_00000_001110; 	// lt
		disk[924] <= 32'b010101_10111_00000_0000001110100111; 	// jf
		disk[925] <= 32'b010001_11101_00111_0000000001100000; 	// la
		disk[926] <= 32'b000000_00111_00101_01111_00000_000000; 	// add
		disk[927] <= 32'b001111_01111_01111_0000000000000000; 	// lw
		disk[928] <= 32'b000010_00101_10000_0000000000000001; 	// subi
		disk[929] <= 32'b000000_00111_10000_10001_00000_000000; 	// add
		disk[930] <= 32'b010010_10001_01111_0000000000000000; 	// sw
		disk[931] <= 32'b000001_00101_10010_0000000000000001; 	// addi
		disk[932] <= 32'b010010_11110_10010_0000000000000000; 	// sw
		disk[933] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[934] <= 32'b111100_00000000000000001110011001; 	// j
		disk[935] <= 32'b001111_11101_00101_0000000011101110; 	// lw
		disk[936] <= 32'b000010_00101_10011_0000000000000001; 	// subi
		disk[937] <= 32'b010001_11101_00110_0000000001100000; 	// la
		disk[938] <= 32'b000000_00110_10011_10100_00000_000000; 	// add
		disk[939] <= 32'b010000_00000_10101_0000000000000000; 	// li
		disk[940] <= 32'b010010_10100_10101_0000000000000000; 	// sw
		disk[941] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[942] <= 32'b000001_11110_11110_0000000000000011; 	// addi
		disk[943] <= 32'b010000_00000_01111_0000000000000001; 	// li
		disk[944] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[945] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[946] <= 32'b001111_11101_00110_0000000011101110; 	// lw
		disk[947] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
		disk[948] <= 32'b010101_10000_00000_0000001110111111; 	// jf
		disk[949] <= 32'b010001_11101_00111_0000000001100000; 	// la
		disk[950] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
		disk[951] <= 32'b001111_10001_10001_0000000000000000; 	// lw
		disk[952] <= 32'b000010_00101_10010_0000000000000001; 	// subi
		disk[953] <= 32'b000000_00111_10010_10011_00000_000000; 	// add
		disk[954] <= 32'b010010_10011_10001_0000000000000000; 	// sw
		disk[955] <= 32'b000001_00101_10100_0000000000000001; 	// addi
		disk[956] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[957] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[958] <= 32'b111100_00000000000000001110110001; 	// j
		disk[959] <= 32'b001111_11101_00101_0000000011101110; 	// lw
		disk[960] <= 32'b000010_00101_10101_0000000000000001; 	// subi
		disk[961] <= 32'b010001_11101_00110_0000000001100000; 	// la
		disk[962] <= 32'b000000_00110_10101_10110_00000_000000; 	// add
		disk[963] <= 32'b010000_00000_10111_0000000000000000; 	// li
		disk[964] <= 32'b010010_10110_10111_0000000000000000; 	// sw
		disk[965] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[966] <= 32'b000001_11110_11110_0000000000000011; 	// addi
		disk[967] <= 32'b010001_11101_00101_0000000001100000; 	// la
		disk[968] <= 32'b001111_00101_01111_0000000000000000; 	// lw
		disk[969] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[970] <= 32'b000000_01111_10001_10000_00000_001101; 	// ne
		disk[971] <= 32'b010101_10000_00000_0000001111010110; 	// jf
		disk[972] <= 32'b001111_00101_10010_0000000000000000; 	// lw
		disk[973] <= 32'b010010_11110_10010_0000000000000000; 	// sw
		disk[974] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[975] <= 32'b111110_00000000000000001110101110; 	// jal
		disk[976] <= 32'b000010_11110_11110_0000000000000011; 	// subi
		disk[977] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[978] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[979] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[980] <= 32'b001110_00110_11000_0000000000000000; 	// mov
		disk[981] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[982] <= 32'b001111_11101_00101_0000000000000011; 	// lw
		disk[983] <= 32'b001110_00101_11000_0000000000000000; 	// mov
		disk[984] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[985] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[986] <= 32'b010010_11110_00001_1111111111111111; 	// sw
		disk[987] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[988] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[989] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[990] <= 32'b001111_11101_00110_0000000011101110; 	// lw
		disk[991] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
		disk[992] <= 32'b010101_10000_00000_0000001111110000; 	// jf
		disk[993] <= 32'b010001_11101_00111_0000000001100000; 	// la
		disk[994] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
		disk[995] <= 32'b001111_10001_10001_0000000000000000; 	// lw
		disk[996] <= 32'b010000_00000_10011_0000000000000000; 	// li
		disk[997] <= 32'b000000_10001_10011_10010_00000_001100; 	// eq
		disk[998] <= 32'b010101_10010_00000_0000001111101011; 	// jf
		disk[999] <= 32'b000000_00111_00101_10100_00000_000000; 	// add
		disk[1000] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[1001] <= 32'b010010_10100_01000_0000000000000000; 	// sw
		disk[1002] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1003] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1004] <= 32'b000001_00101_10101_0000000000000001; 	// addi
		disk[1005] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[1006] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1007] <= 32'b111100_00000000000000001111011101; 	// j
		disk[1008] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1009] <= 32'b000001_11110_11110_0000000000000011; 	// addi
		disk[1010] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[1011] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[1012] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1013] <= 32'b001111_11101_00110_0000000011101110; 	// lw
		disk[1014] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
		disk[1015] <= 32'b010101_10000_00000_0000010000010011; 	// jf
		disk[1016] <= 32'b010001_11101_00111_0000000110010100; 	// la
		disk[1017] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
		disk[1018] <= 32'b001111_10001_10001_0000000000000000; 	// lw
		disk[1019] <= 32'b010000_00000_10011_0000000000000000; 	// li
		disk[1020] <= 32'b000000_10001_10011_10010_00000_001101; 	// ne
		disk[1021] <= 32'b010101_10010_00000_0000010000001110; 	// jf
		disk[1022] <= 32'b010001_11101_01000_0000000000000100; 	// la
		disk[1023] <= 32'b000000_01000_00101_10100_00000_000000; 	// add
		disk[1024] <= 32'b001111_10100_10100_0000000000000000; 	// lw
		disk[1025] <= 32'b001111_11101_01001_0000000000000010; 	// lw
		disk[1026] <= 32'b000000_10100_01001_10101_00000_001101; 	// ne
		disk[1027] <= 32'b010101_10101_00000_0000010000001110; 	// jf
		disk[1028] <= 32'b000000_01000_00101_10110_00000_000000; 	// add
		disk[1029] <= 32'b001111_11101_01010_0000000000000001; 	// lw
		disk[1030] <= 32'b010010_10110_01010_0000000000000000; 	// sw
		disk[1031] <= 32'b000001_00101_10111_0000000000000001; 	// addi
		disk[1032] <= 32'b001110_10111_00001_0000000000000000; 	// mov
		disk[1033] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1034] <= 32'b111110_00000000000000001111011001; 	// jal
		disk[1035] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[1036] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1037] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1038] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1039] <= 32'b000001_00101_01111_0000000000000001; 	// addi
		disk[1040] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[1041] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1042] <= 32'b111100_00000000000000001111110100; 	// j
		disk[1043] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1044] <= 32'b000001_11110_11110_0000000000000101; 	// addi
		disk[1045] <= 32'b010010_11110_00001_1111111111111110; 	// sw
		disk[1046] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[1047] <= 32'b010010_11110_00101_0000000000000000; 	// sw
		disk[1048] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[1049] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[1050] <= 32'b010110_00001_01111_0000000000000000; 	// ldk
		disk[1051] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[1052] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1053] <= 32'b001101_00101_10000_0000000000011010; 	// srli
		disk[1054] <= 32'b001111_11101_00110_0000000110101000; 	// lw
		disk[1055] <= 32'b000000_10000_00110_10001_00000_001101; 	// ne
		disk[1056] <= 32'b010101_10001_00000_0000010000101010; 	// jf
		disk[1057] <= 32'b001111_11110_00111_0000000000000000; 	// lw
		disk[1058] <= 32'b000001_00111_10010_0000000000000001; 	// addi
		disk[1059] <= 32'b010010_11110_10010_0000000000000000; 	// sw
		disk[1060] <= 32'b001111_11110_00111_0000000000000000; 	// lw
		disk[1061] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[1062] <= 32'b010110_00001_10011_0000000000000000; 	// ldk
		disk[1063] <= 32'b010010_11110_10011_1111111111111111; 	// sw
		disk[1064] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1065] <= 32'b111100_00000000000000010000011100; 	// j
		disk[1066] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1067] <= 32'b001111_11110_00110_1111111111111110; 	// lw
		disk[1068] <= 32'b000000_00101_00110_10100_00000_000001; 	// sub
		disk[1069] <= 32'b001110_10100_11000_0000000000000000; 	// mov
		disk[1070] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1071] <= 32'b000001_11110_11110_0000000000001010; 	// addi
		disk[1072] <= 32'b010010_11110_00001_1111111111111001; 	// sw
		disk[1073] <= 32'b001111_11110_00101_1111111111111001; 	// lw
		disk[1074] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1075] <= 32'b010010_11110_11111_1111111111111000; 	// sw
		disk[1076] <= 32'b111110_00000000000000000010000110; 	// jal
		disk[1077] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[1078] <= 32'b001111_11110_11111_1111111111111000; 	// lw
		disk[1079] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1080] <= 32'b010010_11110_00101_1111111111111001; 	// sw
		disk[1081] <= 32'b001111_11110_00110_1111111111111001; 	// lw
		disk[1082] <= 32'b010010_11101_00110_0000000001011111; 	// sw
		disk[1083] <= 32'b010001_11101_00111_0000000110000000; 	// la
		disk[1084] <= 32'b000000_00111_00110_01111_00000_000000; 	// add
		disk[1085] <= 32'b001111_01111_01111_0000000000000000; 	// lw
		disk[1086] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[1087] <= 32'b010001_11101_01000_0000000101110110; 	// la
		disk[1088] <= 32'b000000_01000_00110_10000_00000_000000; 	// add
		disk[1089] <= 32'b001111_10000_10000_0000000000000000; 	// lw
		disk[1090] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[1091] <= 32'b001111_11110_01001_1111111111111111; 	// lw
		disk[1092] <= 32'b010010_11110_01001_1111111111111010; 	// sw
		disk[1093] <= 32'b001110_01001_00001_0000000000000000; 	// mov
		disk[1094] <= 32'b010010_11110_11111_1111111111111000; 	// sw
		disk[1095] <= 32'b111110_00000000000000010000010100; 	// jal
		disk[1096] <= 32'b000010_11110_11110_0000000000000101; 	// subi
		disk[1097] <= 32'b001111_11110_11111_1111111111111000; 	// lw
		disk[1098] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1099] <= 32'b010010_11110_00101_1111111111111110; 	// sw
		disk[1100] <= 32'b001111_11110_00110_1111111111111110; 	// lw
		disk[1101] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[1102] <= 32'b010010_11110_11111_1111111111111000; 	// sw
		disk[1103] <= 32'b111110_00000000000000001011110011; 	// jal
		disk[1104] <= 32'b000010_11110_11110_0000000000000110; 	// subi
		disk[1105] <= 32'b001111_11110_11111_1111111111111000; 	// lw
		disk[1106] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1107] <= 32'b010010_11110_00101_1111111111111101; 	// sw
		disk[1108] <= 32'b010001_11101_00110_0000000000110110; 	// la
		disk[1109] <= 32'b001111_11101_00111_0000000001011111; 	// lw
		disk[1110] <= 32'b000000_00110_00111_10001_00000_000000; 	// add
		disk[1111] <= 32'b001111_11110_01000_1111111111111101; 	// lw
		disk[1112] <= 32'b010010_10001_01000_0000000000000000; 	// sw
		disk[1113] <= 32'b001111_11101_01001_0000000011101011; 	// lw
		disk[1114] <= 32'b000000_01001_01000_10010_00000_000010; 	// mul
		disk[1115] <= 32'b010010_11110_10010_1111111111111011; 	// sw
		disk[1116] <= 32'b001111_11110_01010_1111111111111010; 	// lw
		disk[1117] <= 32'b001110_01010_00001_0000000000000000; 	// mov
		disk[1118] <= 32'b010110_00001_10011_0000000000000000; 	// ldk
		disk[1119] <= 32'b010010_11110_10011_1111111111111100; 	// sw
		disk[1120] <= 32'b001111_11110_00101_1111111111111100; 	// lw
		disk[1121] <= 32'b001101_00101_10100_0000000000011010; 	// srli
		disk[1122] <= 32'b001111_11101_00110_0000000110101000; 	// lw
		disk[1123] <= 32'b000000_10100_00110_10101_00000_001101; 	// ne
		disk[1124] <= 32'b010101_10101_00000_0000010001110101; 	// jf
		disk[1125] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1126] <= 32'b001111_11110_00111_1111111111111011; 	// lw
		disk[1127] <= 32'b001110_00111_00010_0000000000000000; 	// mov
		disk[1128] <= 32'b011001_00010_00001_0000000000000000; 	// sim
		disk[1129] <= 32'b001111_11110_01000_1111111111111010; 	// lw
		disk[1130] <= 32'b000001_01000_10110_0000000000000001; 	// addi
		disk[1131] <= 32'b010010_11110_10110_1111111111111010; 	// sw
		disk[1132] <= 32'b001111_11110_01000_1111111111111010; 	// lw
		disk[1133] <= 32'b001110_01000_00001_0000000000000000; 	// mov
		disk[1134] <= 32'b010110_00001_10111_0000000000000000; 	// ldk
		disk[1135] <= 32'b010010_11110_10111_1111111111111100; 	// sw
		disk[1136] <= 32'b001111_11110_00101_1111111111111100; 	// lw
		disk[1137] <= 32'b000001_00111_01111_0000000000000001; 	// addi
		disk[1138] <= 32'b010010_11110_01111_1111111111111011; 	// sw
		disk[1139] <= 32'b001111_11110_00111_1111111111111011; 	// lw
		disk[1140] <= 32'b111100_00000000000000010001100000; 	// j
		disk[1141] <= 32'b001111_11110_00101_1111111111111100; 	// lw
		disk[1142] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1143] <= 32'b001111_11110_00110_1111111111111011; 	// lw
		disk[1144] <= 32'b001110_00110_00010_0000000000000000; 	// mov
		disk[1145] <= 32'b011001_00010_00001_0000000000000000; 	// sim
		disk[1146] <= 32'b001111_11110_00111_0000000000000000; 	// lw
		disk[1147] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[1148] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
		disk[1149] <= 32'b001111_11101_01000_0000000011101011; 	// lw
		disk[1150] <= 32'b001111_11110_01001_1111111111111101; 	// lw
		disk[1151] <= 32'b000000_01000_01001_10000_00000_000010; 	// mul
		disk[1152] <= 32'b001110_10000_00001_0000000000000000; 	// mov
		disk[1153] <= 32'b011010_00000_00001_0000000000000000; 	// mmuLowerIM
		disk[1154] <= 32'b010001_11101_01010_0000000110010100; 	// la
		disk[1155] <= 32'b001111_11110_01011_1111111111111001; 	// lw
		disk[1156] <= 32'b000000_01010_01011_10001_00000_000000; 	// add
		disk[1157] <= 32'b010010_10001_00111_0000000000000000; 	// sw
		disk[1158] <= 32'b010001_11101_01100_0000000110011110; 	// la
		disk[1159] <= 32'b000000_01100_01011_10010_00000_000000; 	// add
		disk[1160] <= 32'b001111_11110_01101_1111111111111111; 	// lw
		disk[1161] <= 32'b010010_10010_01101_0000000000000000; 	// sw
		disk[1162] <= 32'b010000_00000_10011_0000000000000000; 	// li
		disk[1163] <= 32'b010010_11101_10011_0000000001011111; 	// sw
		disk[1164] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1165] <= 32'b000001_11110_11110_0000000000000110; 	// addi
		disk[1166] <= 32'b001111_11101_00101_0000000011101111; 	// lw
		disk[1167] <= 32'b010010_11110_00101_1111111111111110; 	// sw
		disk[1168] <= 32'b001111_11101_00110_0000000110110000; 	// lw
		disk[1169] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[1170] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[1171] <= 32'b010011_00000_01111_0000000000000000; 	// in
		disk[1172] <= 32'b010010_11110_01111_1111111111111101; 	// sw
		disk[1173] <= 32'b001111_11110_00111_1111111111111101; 	// lw
		disk[1174] <= 32'b000010_00111_10000_0000000000000001; 	// subi
		disk[1175] <= 32'b010010_11110_10000_1111111111111101; 	// sw
		disk[1176] <= 32'b001111_11110_00111_1111111111111101; 	// lw
		disk[1177] <= 32'b000001_00111_10001_0000000000000001; 	// addi
		disk[1178] <= 32'b010001_11101_01000_0000000101110110; 	// la
		disk[1179] <= 32'b000000_01000_00111_10010_00000_000000; 	// add
		disk[1180] <= 32'b010010_10010_10001_0000000000000000; 	// sw
		disk[1181] <= 32'b000000_01000_00111_10011_00000_000000; 	// add
		disk[1182] <= 32'b001111_10011_10011_0000000000000000; 	// lw
		disk[1183] <= 32'b010001_11101_01001_0000000110001010; 	// la
		disk[1184] <= 32'b000000_01001_00111_10100_00000_000000; 	// add
		disk[1185] <= 32'b010010_10100_10011_0000000000000000; 	// sw
		disk[1186] <= 32'b010001_11101_01010_0000000110000000; 	// la
		disk[1187] <= 32'b000000_01010_00111_10101_00000_000000; 	// add
		disk[1188] <= 32'b001111_11110_01011_1111111111111110; 	// lw
		disk[1189] <= 32'b010010_10101_01011_0000000000000000; 	// sw
		disk[1190] <= 32'b001111_11101_01100_0000000110101001; 	// lw
		disk[1191] <= 32'b010010_11110_01100_1111111111111111; 	// sw
		disk[1192] <= 32'b001111_11110_01101_1111111111111111; 	// lw
		disk[1193] <= 32'b001100_01101_10110_0000000000011010; 	// slli
		disk[1194] <= 32'b010010_11110_10110_1111111111111111; 	// sw
		disk[1195] <= 32'b001111_11110_01101_1111111111111111; 	// lw
		disk[1196] <= 32'b000001_01101_10111_0000000000000001; 	// addi
		disk[1197] <= 32'b010010_11110_10111_1111111111111111; 	// sw
		disk[1198] <= 32'b001111_11110_01101_1111111111111111; 	// lw
		disk[1199] <= 32'b001110_01101_00001_0000000000000000; 	// mov
		disk[1200] <= 32'b001110_01011_00010_0000000000000000; 	// mov
		disk[1201] <= 32'b010111_00010_00001_0000000000000000; 	// sdk
		disk[1202] <= 32'b000001_01011_01111_0000000000000001; 	// addi
		disk[1203] <= 32'b010010_11110_01111_1111111111111110; 	// sw
		disk[1204] <= 32'b001111_11110_01011_1111111111111110; 	// lw
		disk[1205] <= 32'b001111_11101_01110_0000000110110001; 	// lw
		disk[1206] <= 32'b001110_01110_00001_0000000000000000; 	// mov
		disk[1207] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[1208] <= 32'b010011_00000_10000_0000000000000000; 	// in
		disk[1209] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[1210] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1211] <= 32'b010000_00000_10010_0000000000000000; 	// li
		disk[1212] <= 32'b000000_00101_10010_10001_00000_001101; 	// ne
		disk[1213] <= 32'b010101_10001_00000_0000010011110000; 	// jf
		disk[1214] <= 32'b001111_11101_00110_0000000110110010; 	// lw
		disk[1215] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[1216] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[1217] <= 32'b010011_00000_10011_0000000000000000; 	// in
		disk[1218] <= 32'b010010_11110_10011_1111111111111111; 	// sw
		disk[1219] <= 32'b001111_11101_00111_0000000110110011; 	// lw
		disk[1220] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[1221] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[1222] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[1223] <= 32'b001100_01000_10100_0000000000001000; 	// slli
		disk[1224] <= 32'b010010_11110_10100_1111111111111111; 	// sw
		disk[1225] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[1226] <= 32'b010011_00000_10101_0000000000000000; 	// in
		disk[1227] <= 32'b000000_01000_10101_10110_00000_000000; 	// add
		disk[1228] <= 32'b010010_11110_10110_1111111111111111; 	// sw
		disk[1229] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[1230] <= 32'b001111_11101_01001_0000000110110100; 	// lw
		disk[1231] <= 32'b001110_01001_00001_0000000000000000; 	// mov
		disk[1232] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[1233] <= 32'b001100_01000_10111_0000000000001000; 	// slli
		disk[1234] <= 32'b010010_11110_10111_1111111111111111; 	// sw
		disk[1235] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[1236] <= 32'b010011_00000_01111_0000000000000000; 	// in
		disk[1237] <= 32'b000000_01000_01111_10000_00000_000000; 	// add
		disk[1238] <= 32'b010010_11110_10000_1111111111111111; 	// sw
		disk[1239] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[1240] <= 32'b001111_11101_01010_0000000110110101; 	// lw
		disk[1241] <= 32'b001110_01010_00001_0000000000000000; 	// mov
		disk[1242] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[1243] <= 32'b001100_01000_10001_0000000000001000; 	// slli
		disk[1244] <= 32'b010010_11110_10001_1111111111111111; 	// sw
		disk[1245] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[1246] <= 32'b010011_00000_10010_0000000000000000; 	// in
		disk[1247] <= 32'b000000_01000_10010_10011_00000_000000; 	// add
		disk[1248] <= 32'b010010_11110_10011_1111111111111111; 	// sw
		disk[1249] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[1250] <= 32'b001110_01000_00001_0000000000000000; 	// mov
		disk[1251] <= 32'b001111_11110_01011_1111111111111110; 	// lw
		disk[1252] <= 32'b001110_01011_00010_0000000000000000; 	// mov
		disk[1253] <= 32'b010111_00010_00001_0000000000000000; 	// sdk
		disk[1254] <= 32'b000001_01011_10100_0000000000000001; 	// addi
		disk[1255] <= 32'b010010_11110_10100_1111111111111110; 	// sw
		disk[1256] <= 32'b001111_11110_01011_1111111111111110; 	// lw
		disk[1257] <= 32'b001111_11101_01100_0000000110110001; 	// lw
		disk[1258] <= 32'b001110_01100_00001_0000000000000000; 	// mov
		disk[1259] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[1260] <= 32'b010011_00000_10101_0000000000000000; 	// in
		disk[1261] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[1262] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1263] <= 32'b111100_00000000000000010010111010; 	// j
		disk[1264] <= 32'b010000_00000_10110_0000000001111111; 	// li
		disk[1265] <= 32'b010010_11110_10110_1111111111111111; 	// sw
		disk[1266] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1267] <= 32'b001100_00101_10111_0000000000001000; 	// slli
		disk[1268] <= 32'b010010_11110_10111_1111111111111111; 	// sw
		disk[1269] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1270] <= 32'b000001_00101_01111_0000000000100000; 	// addi
		disk[1271] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[1272] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1273] <= 32'b001100_00101_10000_0000000000010001; 	// slli
		disk[1274] <= 32'b010010_11110_10000_1111111111111111; 	// sw
		disk[1275] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1276] <= 32'b001101_00101_10001_0000000000000001; 	// srli
		disk[1277] <= 32'b010010_11110_10001_1111111111111111; 	// sw
		disk[1278] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1279] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1280] <= 32'b001111_11110_00110_1111111111111110; 	// lw
		disk[1281] <= 32'b001110_00110_00010_0000000000000000; 	// mov
		disk[1282] <= 32'b010111_00010_00001_0000000000000000; 	// sdk
		disk[1283] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1284] <= 32'b000001_11110_11110_0000000000000011; 	// addi
		disk[1285] <= 32'b010010_11110_00001_0000000000000000; 	// sw
		disk[1286] <= 32'b010001_11101_00101_0000000110010100; 	// la
		disk[1287] <= 32'b001111_11101_00110_0000000001011111; 	// lw
		disk[1288] <= 32'b000000_00101_00110_01111_00000_000000; 	// add
		disk[1289] <= 32'b001111_01111_01111_0000000000000000; 	// lw
		disk[1290] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[1291] <= 32'b000000_01111_10001_10000_00000_001101; 	// ne
		disk[1292] <= 32'b010101_10000_00000_0000010100111000; 	// jf
		disk[1293] <= 32'b001111_11110_00111_0000000000000000; 	// lw
		disk[1294] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[1295] <= 32'b100100_00000_00001_0000000000000000; 	// lcdCurr
		disk[1296] <= 32'b001111_11101_01000_0000000110111100; 	// lw
		disk[1297] <= 32'b001110_01000_00001_0000000000000000; 	// mov
		disk[1298] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[1299] <= 32'b001111_11101_01001_0000000011110001; 	// lw
		disk[1300] <= 32'b000001_01001_10010_0000000000000001; 	// addi
		disk[1301] <= 32'b010010_11101_10010_0000000011110010; 	// sw
		disk[1302] <= 32'b010001_11101_01010_0000000000000100; 	// la
		disk[1303] <= 32'b000000_01010_00110_10011_00000_000000; 	// add
		disk[1304] <= 32'b001111_11101_01011_0000000000000000; 	// lw
		disk[1305] <= 32'b010010_10011_01011_0000000000000000; 	// sw
		disk[1306] <= 32'b010001_11101_01100_0000000000001110; 	// la
		disk[1307] <= 32'b000000_01100_00110_10100_00000_000000; 	// add
		disk[1308] <= 32'b010000_00000_10101_0000000000000000; 	// li
		disk[1309] <= 32'b010010_10100_10101_0000000000000000; 	// sw
		disk[1310] <= 32'b001111_11101_01101_0000000011110010; 	// lw
		disk[1311] <= 32'b001110_01101_00001_0000000000000000; 	// mov
		disk[1312] <= 32'b001110_00001_11100_0000000000000000; 	// mov
		disk[1313] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[1314] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
		disk[1315] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1316] <= 32'b001110_11110_00011_0000000000000000; 	// mov
		disk[1317] <= 32'b001110_11101_00100_0000000000000000; 	// mov
		disk[1318] <= 32'b001110_11100_11110_0000000000000000; 	// mov
		disk[1319] <= 32'b001110_11011_11101_0000000000000000; 	// mov
		disk[1320] <= 32'b001110_00011_11100_0000000000000000; 	// mov
		disk[1321] <= 32'b001110_00100_11011_0000000000000000; 	// mov
		disk[1322] <= 32'b100000_00000000000000000000000000; 	// exec
		disk[1323] <= 32'b001110_11100_11110_0000000000000000; 	// mov
		disk[1324] <= 32'b001110_11011_11101_0000000000000000; 	// mov
		disk[1325] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1326] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1327] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1328] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1329] <= 32'b111110_00000000000000000010100000; 	// jal
		disk[1330] <= 32'b000010_11110_11110_0000000000000101; 	// subi
		disk[1331] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1332] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1333] <= 32'b001111_11101_00110_0000000110101011; 	// lw
		disk[1334] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[1335] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[1336] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1337] <= 32'b000001_11110_11110_0000000000001000; 	// addi
		disk[1338] <= 32'b010010_11110_00001_1111111111111011; 	// sw
		disk[1339] <= 32'b001111_11110_00101_1111111111111011; 	// lw
		disk[1340] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1341] <= 32'b100100_00000_00001_0000000000000000; 	// lcdCurr
		disk[1342] <= 32'b001111_11101_00110_0000000110111100; 	// lw
		disk[1343] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[1344] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[1345] <= 32'b001111_11101_00111_0000000011110001; 	// lw
		disk[1346] <= 32'b000001_00111_01111_0000000000000001; 	// addi
		disk[1347] <= 32'b010010_11101_01111_0000000011110010; 	// sw
		disk[1348] <= 32'b010001_11101_01000_0000000000000100; 	// la
		disk[1349] <= 32'b001111_11101_01001_0000000001011111; 	// lw
		disk[1350] <= 32'b000000_01000_01001_10000_00000_000000; 	// add
		disk[1351] <= 32'b001111_11101_01010_0000000000000000; 	// lw
		disk[1352] <= 32'b010010_10000_01010_0000000000000000; 	// sw
		disk[1353] <= 32'b010001_11101_01011_0000000001000000; 	// la
		disk[1354] <= 32'b000000_01011_01001_10001_00000_000000; 	// add
		disk[1355] <= 32'b001111_10001_10001_0000000000000000; 	// lw
		disk[1356] <= 32'b010010_11110_10001_1111111111111101; 	// sw
		disk[1357] <= 32'b001111_11101_01100_0000000011110010; 	// lw
		disk[1358] <= 32'b010010_11110_01100_1111111111111110; 	// sw
		disk[1359] <= 32'b001111_11110_01101_1111111111111101; 	// lw
		disk[1360] <= 32'b001111_11101_01110_0000000011101011; 	// lw
		disk[1361] <= 32'b000000_01101_01110_10010_00000_000010; 	// mul
		disk[1362] <= 32'b010010_11110_10010_1111111111111111; 	// sw
		disk[1363] <= 32'b010001_11101_00101_0000000000011000; 	// la
		disk[1364] <= 32'b000000_00101_01001_10011_00000_000000; 	// add
		disk[1365] <= 32'b001111_10011_10011_0000000000000000; 	// lw
		disk[1366] <= 32'b010010_11110_10011_0000000000000000; 	// sw
		disk[1367] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1368] <= 32'b010000_00000_10101_0000000000000000; 	// li
		disk[1369] <= 32'b000000_00101_10101_10100_00000_010000; 	// gt
		disk[1370] <= 32'b010101_10100_00000_0000010101101110; 	// jf
		disk[1371] <= 32'b001111_11110_00110_1111111111111111; 	// lw
		disk[1372] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[1373] <= 32'b001111_00001_10110_0000000000000000; 	// lw
		disk[1374] <= 32'b010010_11110_10110_1111111111111100; 	// sw
		disk[1375] <= 32'b001111_11110_00111_1111111111111100; 	// lw
		disk[1376] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[1377] <= 32'b001111_11110_01000_1111111111111110; 	// lw
		disk[1378] <= 32'b001110_01000_00010_0000000000000000; 	// mov
		disk[1379] <= 32'b010010_00010_00001_0000000000000000; 	// sw
		disk[1380] <= 32'b000001_01000_10111_0000000000000001; 	// addi
		disk[1381] <= 32'b010010_11110_10111_1111111111111110; 	// sw
		disk[1382] <= 32'b001111_11110_01000_1111111111111110; 	// lw
		disk[1383] <= 32'b000001_00110_01111_0000000000000001; 	// addi
		disk[1384] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[1385] <= 32'b001111_11110_00110_1111111111111111; 	// lw
		disk[1386] <= 32'b000010_00101_10000_0000000000000001; 	// subi
		disk[1387] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[1388] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1389] <= 32'b111100_00000000000000010101010111; 	// j
		disk[1390] <= 32'b010001_11101_00101_0000000000011000; 	// la
		disk[1391] <= 32'b001111_11101_00110_0000000001011111; 	// lw
		disk[1392] <= 32'b000000_00101_00110_10001_00000_000000; 	// add
		disk[1393] <= 32'b001111_10001_10001_0000000000000000; 	// lw
		disk[1394] <= 32'b001111_11101_00111_0000000011110001; 	// lw
		disk[1395] <= 32'b000000_00111_10001_10010_00000_000000; 	// add
		disk[1396] <= 32'b001110_10010_00001_0000000000000000; 	// mov
		disk[1397] <= 32'b001110_00001_11100_0000000000000000; 	// mov
		disk[1398] <= 32'b000001_00110_10011_0000000000000001; 	// addi
		disk[1399] <= 32'b001110_10011_00001_0000000000000000; 	// mov
		disk[1400] <= 32'b010001_11101_01000_0000000000001110; 	// la
		disk[1401] <= 32'b000000_01000_00110_10100_00000_000000; 	// add
		disk[1402] <= 32'b001111_10100_10100_0000000000000000; 	// lw
		disk[1403] <= 32'b001110_10100_00010_0000000000000000; 	// mov
		disk[1404] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
		disk[1405] <= 32'b010010_11110_11111_1111111111111010; 	// sw
		disk[1406] <= 32'b001110_11110_00011_0000000000000000; 	// mov
		disk[1407] <= 32'b001110_11101_00100_0000000000000000; 	// mov
		disk[1408] <= 32'b001110_11100_11110_0000000000000000; 	// mov
		disk[1409] <= 32'b001110_11011_11101_0000000000000000; 	// mov
		disk[1410] <= 32'b001110_00011_11100_0000000000000000; 	// mov
		disk[1411] <= 32'b001110_00100_11011_0000000000000000; 	// mov
		disk[1412] <= 32'b001110_00010_11010_0000000000000000; 	// mov
		disk[1413] <= 32'b001111_00000_00000_0000111111100000; 	// lw
		disk[1414] <= 32'b001111_00000_00001_0000111111100001; 	// lw
		disk[1415] <= 32'b001111_00000_00010_0000111111100010; 	// lw
		disk[1416] <= 32'b001111_00000_00011_0000111111100011; 	// lw
		disk[1417] <= 32'b001111_00000_00100_0000111111100100; 	// lw
		disk[1418] <= 32'b001111_00000_00101_0000111111100101; 	// lw
		disk[1419] <= 32'b001111_00000_00110_0000111111100110; 	// lw
		disk[1420] <= 32'b001111_00000_00111_0000111111100111; 	// lw
		disk[1421] <= 32'b001111_00000_01000_0000111111101000; 	// lw
		disk[1422] <= 32'b001111_00000_01001_0000111111101001; 	// lw
		disk[1423] <= 32'b001111_00000_01010_0000111111101010; 	// lw
		disk[1424] <= 32'b001111_00000_01011_0000111111101011; 	// lw
		disk[1425] <= 32'b001111_00000_01100_0000111111101100; 	// lw
		disk[1426] <= 32'b001111_00000_01101_0000111111101101; 	// lw
		disk[1427] <= 32'b001111_00000_01110_0000111111101110; 	// lw
		disk[1428] <= 32'b001111_00000_01111_0000111111101111; 	// lw
		disk[1429] <= 32'b001111_00000_10000_0000111111110000; 	// lw
		disk[1430] <= 32'b001111_00000_10001_0000111111110001; 	// lw
		disk[1431] <= 32'b001111_00000_10010_0000111111110010; 	// lw
		disk[1432] <= 32'b001111_00000_10011_0000111111110011; 	// lw
		disk[1433] <= 32'b001111_00000_10100_0000111111110100; 	// lw
		disk[1434] <= 32'b001111_00000_10101_0000111111110101; 	// lw
		disk[1435] <= 32'b001111_00000_10110_0000111111110110; 	// lw
		disk[1436] <= 32'b001111_00000_10111_0000111111110111; 	// lw
		disk[1437] <= 32'b001111_00000_11000_0000111111111000; 	// lw
		disk[1438] <= 32'b001111_00000_11111_0000111111111001; 	// lw
		disk[1439] <= 32'b100001_11010_00000_0000000000000000; 	// execAgain
		disk[1440] <= 32'b001110_11100_11110_0000000000000000; 	// mov
		disk[1441] <= 32'b001110_11011_11101_0000000000000000; 	// mov
		disk[1442] <= 32'b001111_11110_11111_1111111111111010; 	// lw
		disk[1443] <= 32'b001111_11110_00101_1111111111111011; 	// lw
		disk[1444] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1445] <= 32'b010010_11110_11111_1111111111111010; 	// sw
		disk[1446] <= 32'b111110_00000000000000000010100000; 	// jal
		disk[1447] <= 32'b000010_11110_11110_0000000000000101; 	// subi
		disk[1448] <= 32'b001111_11110_11111_1111111111111010; 	// lw
		disk[1449] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1450] <= 32'b001111_11101_00110_0000000110101011; 	// lw
		disk[1451] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[1452] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[1453] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1454] <= 32'b000001_11110_11110_0000000000000011; 	// addi
		disk[1455] <= 32'b010010_11110_00001_0000000000000000; 	// sw
		disk[1456] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1457] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1458] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1459] <= 32'b111110_00000000000000000010000110; 	// jal
		disk[1460] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[1461] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1462] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1463] <= 32'b010010_11101_00101_0000000001011111; 	// sw
		disk[1464] <= 32'b001111_11101_00110_0000000001011111; 	// lw
		disk[1465] <= 32'b000001_00110_01111_0000000000000001; 	// addi
		disk[1466] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[1467] <= 32'b010010_11101_00110_0000000001011110; 	// sw
		disk[1468] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1469] <= 32'b111110_00000000000000000000111110; 	// jal
		disk[1470] <= 32'b000010_11110_11110_0000000000000110; 	// subi
		disk[1471] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1472] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1473] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[1474] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[1475] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1476] <= 32'b111110_00000000000000010100111001; 	// jal
		disk[1477] <= 32'b000010_11110_11110_0000000000001000; 	// subi
		disk[1478] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1479] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1480] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1481] <= 32'b000001_11110_11110_0000000000000011; 	// addi
		disk[1482] <= 32'b010010_11110_00001_0000000000000000; 	// sw
		disk[1483] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1484] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1485] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1486] <= 32'b111110_00000000000000000010000110; 	// jal
		disk[1487] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[1488] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1489] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1490] <= 32'b010010_11101_00101_0000000001011111; 	// sw
		disk[1491] <= 32'b001111_11101_00110_0000000001011111; 	// lw
		disk[1492] <= 32'b000001_00110_01111_0000000000000001; 	// addi
		disk[1493] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[1494] <= 32'b010010_11101_00110_0000000001011110; 	// sw
		disk[1495] <= 32'b001111_11110_00111_0000000000000000; 	// lw
		disk[1496] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[1497] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1498] <= 32'b111110_00000000000000010100000100; 	// jal
		disk[1499] <= 32'b000010_11110_11110_0000000000000011; 	// subi
		disk[1500] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1501] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1502] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1503] <= 32'b000001_11110_11110_0000000000000011; 	// addi
		disk[1504] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1505] <= 32'b111110_00000000000000001111110001; 	// jal
		disk[1506] <= 32'b000010_11110_11110_0000000000000011; 	// subi
		disk[1507] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1508] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1509] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1510] <= 32'b111110_00000000000000001111000110; 	// jal
		disk[1511] <= 32'b000010_11110_11110_0000000000000011; 	// subi
		disk[1512] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1513] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1514] <= 32'b010010_11110_00101_0000000000000000; 	// sw
		disk[1515] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1516] <= 32'b001111_11101_00110_0000000000000011; 	// lw
		disk[1517] <= 32'b000000_00101_00110_01111_00000_001101; 	// ne
		disk[1518] <= 32'b010101_01111_00000_0000011000010010; 	// jf
		disk[1519] <= 32'b000010_00101_10000_0000000000000001; 	// subi
		disk[1520] <= 32'b010010_11101_10000_0000000001011111; 	// sw
		disk[1521] <= 32'b010001_11101_00111_0000000000001110; 	// la
		disk[1522] <= 32'b001111_11101_01000_0000000001011111; 	// lw
		disk[1523] <= 32'b000000_00111_01000_10001_00000_000000; 	// add
		disk[1524] <= 32'b001111_10001_10001_0000000000000000; 	// lw
		disk[1525] <= 32'b010000_00000_10011_0000000000000000; 	// li
		disk[1526] <= 32'b000000_10001_10011_10010_00000_001100; 	// eq
		disk[1527] <= 32'b010101_10010_00000_0000010111111111; 	// jf
		disk[1528] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1529] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1530] <= 32'b111110_00000000000000010100000100; 	// jal
		disk[1531] <= 32'b000010_11110_11110_0000000000000011; 	// subi
		disk[1532] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1533] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1534] <= 32'b111100_00000000000000011000001011; 	// j
		disk[1535] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1536] <= 32'b111110_00000000000000000000111110; 	// jal
		disk[1537] <= 32'b000010_11110_11110_0000000000000110; 	// subi
		disk[1538] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1539] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1540] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[1541] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[1542] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1543] <= 32'b111110_00000000000000010100111001; 	// jal
		disk[1544] <= 32'b000010_11110_11110_0000000000001000; 	// subi
		disk[1545] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1546] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1547] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1548] <= 32'b111110_00000000000000001111000110; 	// jal
		disk[1549] <= 32'b000010_11110_11110_0000000000000011; 	// subi
		disk[1550] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1551] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1552] <= 32'b010010_11110_00101_0000000000000000; 	// sw
		disk[1553] <= 32'b111100_00000000000000010111101011; 	// j
		disk[1554] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[1555] <= 32'b010010_11101_10100_0000000001101010; 	// sw
		disk[1556] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1557] <= 32'b001110_11110_11100_0000000000000000; 	// mov
		disk[1558] <= 32'b001110_11101_11011_0000000000000000; 	// mov
		disk[1559] <= 32'b010000_00000_00000_0000000000000000; 	// li
		disk[1560] <= 32'b010000_00000_11110_0000000000000000; 	// li
		disk[1561] <= 32'b010000_00000_11101_0000000000000000; 	// li
		disk[1562] <= 32'b000001_11110_11110_0000000111000111; 	// addi
		disk[1563] <= 32'b010010_00000_00000_0000111111100000; 	// sw
		disk[1564] <= 32'b010010_00000_00001_0000111111100001; 	// sw
		disk[1565] <= 32'b010010_00000_00010_0000111111100010; 	// sw
		disk[1566] <= 32'b010010_00000_00011_0000111111100011; 	// sw
		disk[1567] <= 32'b010010_00000_00100_0000111111100100; 	// sw
		disk[1568] <= 32'b010010_00000_00101_0000111111100101; 	// sw
		disk[1569] <= 32'b010010_00000_00110_0000111111100110; 	// sw
		disk[1570] <= 32'b010010_00000_00111_0000111111100111; 	// sw
		disk[1571] <= 32'b010010_00000_01000_0000111111101000; 	// sw
		disk[1572] <= 32'b010010_00000_01001_0000111111101001; 	// sw
		disk[1573] <= 32'b010010_00000_01010_0000111111101010; 	// sw
		disk[1574] <= 32'b010010_00000_01011_0000111111101011; 	// sw
		disk[1575] <= 32'b010010_00000_01100_0000111111101100; 	// sw
		disk[1576] <= 32'b010010_00000_01101_0000111111101101; 	// sw
		disk[1577] <= 32'b010010_00000_01110_0000111111101110; 	// sw
		disk[1578] <= 32'b010010_00000_01111_0000111111101111; 	// sw
		disk[1579] <= 32'b010010_00000_10000_0000111111110000; 	// sw
		disk[1580] <= 32'b010010_00000_10001_0000111111110001; 	// sw
		disk[1581] <= 32'b010010_00000_10010_0000111111110010; 	// sw
		disk[1582] <= 32'b010010_00000_10011_0000111111110011; 	// sw
		disk[1583] <= 32'b010010_00000_10100_0000111111110100; 	// sw
		disk[1584] <= 32'b010010_00000_10101_0000111111110101; 	// sw
		disk[1585] <= 32'b010010_00000_10110_0000111111110110; 	// sw
		disk[1586] <= 32'b010010_00000_10111_0000111111110111; 	// sw
		disk[1587] <= 32'b010010_00000_11000_0000111111111000; 	// sw
		disk[1588] <= 32'b010010_00000_11111_0000111111111001; 	// sw
		disk[1589] <= 32'b001111_11110_00101_1111111111111011; 	// lw
		disk[1590] <= 32'b010000_00000_10000_0000000000000000; 	// li
		disk[1591] <= 32'b000000_00101_10000_01111_00000_001100; 	// eq
		disk[1592] <= 32'b010101_01111_00000_0000011001000010; 	// jf
		disk[1593] <= 32'b111110_00000000000000001011001110; 	// jal
		disk[1594] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[1595] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1596] <= 32'b001111_11101_00110_0000000110101011; 	// lw
		disk[1597] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[1598] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[1599] <= 32'b010000_00000_10001_0000000000000001; 	// li
		disk[1600] <= 32'b010010_11110_10001_1111111111111011; 	// sw
		disk[1601] <= 32'b100110_00000_00000_0000000000000000; 	// cic
		disk[1602] <= 32'b100101_00000_10010_0000000000000000; 	// gic
		disk[1603] <= 32'b010010_11110_10010_1111111111111010; 	// sw
		disk[1604] <= 32'b001111_11110_00101_1111111111111010; 	// lw
		disk[1605] <= 32'b001111_11101_00110_0000000101110101; 	// lw
		disk[1606] <= 32'b000000_00101_00110_10011_00000_001100; 	// eq
		disk[1607] <= 32'b010101_10011_00000_0000011010111111; 	// jf
		disk[1608] <= 32'b001110_11100_10100_0000000000000000; 	// mov
		disk[1609] <= 32'b010010_11101_10100_0000000011110011; 	// sw
		disk[1610] <= 32'b001111_11101_00111_0000000011110011; 	// lw
		disk[1611] <= 32'b001111_11101_01000_0000000011110010; 	// lw
		disk[1612] <= 32'b000000_00111_01000_10101_00000_000001; 	// sub
		disk[1613] <= 32'b000001_10101_10110_0000000000000001; 	// addi
		disk[1614] <= 32'b010010_11110_10110_0000000000000000; 	// sw
		disk[1615] <= 32'b010001_11101_01001_0000000000011000; 	// la
		disk[1616] <= 32'b001111_11101_01010_0000000001011111; 	// lw
		disk[1617] <= 32'b000000_01001_01010_10111_00000_000000; 	// add
		disk[1618] <= 32'b001111_11110_01011_0000000000000000; 	// lw
		disk[1619] <= 32'b010010_10111_01011_0000000000000000; 	// sw
		disk[1620] <= 32'b010001_11101_01100_0000000000000100; 	// la
		disk[1621] <= 32'b000000_01100_01010_01111_00000_000000; 	// add
		disk[1622] <= 32'b001111_11101_01101_0000000000000010; 	// lw
		disk[1623] <= 32'b010010_01111_01101_0000000000000000; 	// sw
		disk[1624] <= 32'b100111_00000_10000_0000000000000000; 	// gip
		disk[1625] <= 32'b010001_11101_01110_0000000000001110; 	// la
		disk[1626] <= 32'b000000_01110_01010_10001_00000_000000; 	// add
		disk[1627] <= 32'b010010_10001_10000_0000000000000000; 	// sw
		disk[1628] <= 32'b010001_11101_00101_0000000001000000; 	// la
		disk[1629] <= 32'b000000_00101_01010_10010_00000_000000; 	// add
		disk[1630] <= 32'b001111_10010_10010_0000000000000000; 	// lw
		disk[1631] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[1632] <= 32'b000000_10010_10100_10011_00000_001100; 	// eq
		disk[1633] <= 32'b010101_10011_00000_0000011001101100; 	// jf
		disk[1634] <= 32'b111110_00000000000000001100101110; 	// jal
		disk[1635] <= 32'b000010_11110_11110_0000000000000101; 	// subi
		disk[1636] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1637] <= 32'b010010_11110_00101_1111111111111100; 	// sw
		disk[1638] <= 32'b010001_11101_00110_0000000001000000; 	// la
		disk[1639] <= 32'b001111_11101_00111_0000000001011111; 	// lw
		disk[1640] <= 32'b000000_00110_00111_10101_00000_000000; 	// add
		disk[1641] <= 32'b001111_11110_01000_1111111111111100; 	// lw
		disk[1642] <= 32'b010010_10101_01000_0000000000000000; 	// sw
		disk[1643] <= 32'b111100_00000000000000011001110001; 	// j
		disk[1644] <= 32'b010001_11101_00101_0000000001000000; 	// la
		disk[1645] <= 32'b001111_11101_00110_0000000001011111; 	// lw
		disk[1646] <= 32'b000000_00101_00110_10110_00000_000000; 	// add
		disk[1647] <= 32'b001111_10110_10110_0000000000000000; 	// lw
		disk[1648] <= 32'b010010_11110_10110_1111111111111100; 	// sw
		disk[1649] <= 32'b001111_11101_00101_0000000011110010; 	// lw
		disk[1650] <= 32'b010010_11110_00101_1111111111111110; 	// sw
		disk[1651] <= 32'b001111_11110_00110_1111111111111100; 	// lw
		disk[1652] <= 32'b001111_11101_00111_0000000011101011; 	// lw
		disk[1653] <= 32'b000000_00110_00111_10111_00000_000010; 	// mul
		disk[1654] <= 32'b010010_11110_10111_1111111111111111; 	// sw
		disk[1655] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1656] <= 32'b010000_00000_10000_0000000000000000; 	// li
		disk[1657] <= 32'b000000_00101_10000_01111_00000_010000; 	// gt
		disk[1658] <= 32'b010101_01111_00000_0000011010001110; 	// jf
		disk[1659] <= 32'b001111_11110_00110_1111111111111110; 	// lw
		disk[1660] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[1661] <= 32'b001111_00001_10001_0000000000000000; 	// lw
		disk[1662] <= 32'b010010_11110_10001_1111111111111101; 	// sw
		disk[1663] <= 32'b001111_11110_00111_1111111111111101; 	// lw
		disk[1664] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[1665] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[1666] <= 32'b001110_01000_00010_0000000000000000; 	// mov
		disk[1667] <= 32'b010010_00010_00001_0000000000000000; 	// sw
		disk[1668] <= 32'b000001_00110_10010_0000000000000001; 	// addi
		disk[1669] <= 32'b010010_11110_10010_1111111111111110; 	// sw
		disk[1670] <= 32'b001111_11110_00110_1111111111111110; 	// lw
		disk[1671] <= 32'b000001_01000_10011_0000000000000001; 	// addi
		disk[1672] <= 32'b010010_11110_10011_1111111111111111; 	// sw
		disk[1673] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[1674] <= 32'b000010_00101_10100_0000000000000001; 	// subi
		disk[1675] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[1676] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1677] <= 32'b111100_00000000000000011001110111; 	// j
		disk[1678] <= 32'b001111_11101_00101_0000000001011111; 	// lw
		disk[1679] <= 32'b001111_11101_00110_0000000001011110; 	// lw
		disk[1680] <= 32'b000000_00101_00110_10101_00000_001100; 	// eq
		disk[1681] <= 32'b010101_10101_00000_0000011010011000; 	// jf
		disk[1682] <= 32'b000001_00101_10110_0000000000000001; 	// addi
		disk[1683] <= 32'b001110_10110_00001_0000000000000000; 	// mov
		disk[1684] <= 32'b111110_00000000000000010100111001; 	// jal
		disk[1685] <= 32'b000010_11110_11110_0000000000001000; 	// subi
		disk[1686] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1687] <= 32'b111100_00000000000000011010110110; 	// j
		disk[1688] <= 32'b001111_11110_00101_1111111111111100; 	// lw
		disk[1689] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1690] <= 32'b111110_00000000000000000001100011; 	// jal
		disk[1691] <= 32'b000010_11110_11110_0000000000000110; 	// subi
		disk[1692] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1693] <= 32'b010001_11101_00110_0000000000000100; 	// la
		disk[1694] <= 32'b001111_11101_00111_0000000001011111; 	// lw
		disk[1695] <= 32'b000000_00110_00111_10111_00000_000000; 	// add
		disk[1696] <= 32'b001111_11101_01000_0000000000000010; 	// lw
		disk[1697] <= 32'b010010_10111_01000_0000000000000000; 	// sw
		disk[1698] <= 32'b000001_00111_01111_0000000000000001; 	// addi
		disk[1699] <= 32'b001110_01111_00001_0000000000000000; 	// mov
		disk[1700] <= 32'b111110_00000000000000001110000001; 	// jal
		disk[1701] <= 32'b000010_11110_11110_0000000000000101; 	// subi
		disk[1702] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1703] <= 32'b001111_11101_00110_0000000001101010; 	// lw
		disk[1704] <= 32'b010000_00000_10001_0000000000000001; 	// li
		disk[1705] <= 32'b000000_00110_10001_10000_00000_001100; 	// eq
		disk[1706] <= 32'b010101_10000_00000_0000011010110110; 	// jf
		disk[1707] <= 32'b001111_11101_00111_0000000110101011; 	// lw
		disk[1708] <= 32'b010010_11101_00111_0000000110111101; 	// sw
		disk[1709] <= 32'b001111_11101_01000_0000000110111101; 	// lw
		disk[1710] <= 32'b001110_01000_00001_0000000000000000; 	// mov
		disk[1711] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[1712] <= 32'b010000_00000_11101_0000000000000000; 	// li
		disk[1713] <= 32'b010000_00000_11110_0000000111000111; 	// li
		disk[1714] <= 32'b100110_00000_00000_0000000000000000; 	// cic
		disk[1715] <= 32'b111110_00000000000000010111011111; 	// jal
		disk[1716] <= 32'b000010_11110_11110_0000000000000011; 	// subi
		disk[1717] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1718] <= 32'b001111_11101_00101_0000000110101011; 	// lw
		disk[1719] <= 32'b010010_11101_00101_0000000110111101; 	// sw
		disk[1720] <= 32'b001111_11101_00110_0000000110111101; 	// lw
		disk[1721] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[1722] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[1723] <= 32'b010000_00000_11101_0000000000000000; 	// li
		disk[1724] <= 32'b010000_00000_11110_0000000111000111; 	// li
		disk[1725] <= 32'b100110_00000_00000_0000000000000000; 	// cic
		disk[1726] <= 32'b111100_00000000000000011100101011; 	// j
		disk[1727] <= 32'b001111_11110_00101_1111111111111010; 	// lw
		disk[1728] <= 32'b001111_11101_00110_0000000101110100; 	// lw
		disk[1729] <= 32'b000000_00101_00110_10010_00000_001100; 	// eq
		disk[1730] <= 32'b010101_10010_00000_0000011100101011; 	// jf
		disk[1731] <= 32'b001110_11100_10011_0000000000000000; 	// mov
		disk[1732] <= 32'b010010_11101_10011_0000000011110011; 	// sw
		disk[1733] <= 32'b001111_11101_00111_0000000011110011; 	// lw
		disk[1734] <= 32'b001111_11101_01000_0000000011110010; 	// lw
		disk[1735] <= 32'b000000_00111_01000_10100_00000_000001; 	// sub
		disk[1736] <= 32'b000001_10100_10101_0000000000000001; 	// addi
		disk[1737] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[1738] <= 32'b010001_11101_01001_0000000000011000; 	// la
		disk[1739] <= 32'b001111_11101_01010_0000000001011111; 	// lw
		disk[1740] <= 32'b000000_01001_01010_10110_00000_000000; 	// add
		disk[1741] <= 32'b001111_11110_01011_0000000000000000; 	// lw
		disk[1742] <= 32'b010010_10110_01011_0000000000000000; 	// sw
		disk[1743] <= 32'b010001_11101_01100_0000000000000100; 	// la
		disk[1744] <= 32'b000000_01100_01010_10111_00000_000000; 	// add
		disk[1745] <= 32'b001111_11101_01101_0000000000000010; 	// lw
		disk[1746] <= 32'b010010_10111_01101_0000000000000000; 	// sw
		disk[1747] <= 32'b100111_00000_01111_0000000000000000; 	// gip
		disk[1748] <= 32'b010001_11101_01110_0000000000001110; 	// la
		disk[1749] <= 32'b000000_01110_01010_10000_00000_000000; 	// add
		disk[1750] <= 32'b010010_10000_01111_0000000000000000; 	// sw
		disk[1751] <= 32'b010001_11101_00101_0000000001000000; 	// la
		disk[1752] <= 32'b000000_00101_01010_10001_00000_000000; 	// add
		disk[1753] <= 32'b001111_10001_10001_0000000000000000; 	// lw
		disk[1754] <= 32'b010000_00000_10011_0000000000000000; 	// li
		disk[1755] <= 32'b000000_10001_10011_10010_00000_001100; 	// eq
		disk[1756] <= 32'b010101_10010_00000_0000011011100111; 	// jf
		disk[1757] <= 32'b111110_00000000000000001100101110; 	// jal
		disk[1758] <= 32'b000010_11110_11110_0000000000000101; 	// subi
		disk[1759] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1760] <= 32'b010010_11110_00101_1111111111111100; 	// sw
		disk[1761] <= 32'b010001_11101_00110_0000000001000000; 	// la
		disk[1762] <= 32'b001111_11101_00111_0000000001011111; 	// lw
		disk[1763] <= 32'b000000_00110_00111_10100_00000_000000; 	// add
		disk[1764] <= 32'b001111_11110_01000_1111111111111100; 	// lw
		disk[1765] <= 32'b010010_10100_01000_0000000000000000; 	// sw
		disk[1766] <= 32'b111100_00000000000000011011101100; 	// j
		disk[1767] <= 32'b010001_11101_00101_0000000001000000; 	// la
		disk[1768] <= 32'b001111_11101_00110_0000000001011111; 	// lw
		disk[1769] <= 32'b000000_00101_00110_10101_00000_000000; 	// add
		disk[1770] <= 32'b001111_10101_10101_0000000000000000; 	// lw
		disk[1771] <= 32'b010010_11110_10101_1111111111111100; 	// sw
		disk[1772] <= 32'b001111_11101_00101_0000000011110010; 	// lw
		disk[1773] <= 32'b010010_11110_00101_1111111111111110; 	// sw
		disk[1774] <= 32'b001111_11110_00110_1111111111111100; 	// lw
		disk[1775] <= 32'b001111_11101_00111_0000000011101011; 	// lw
		disk[1776] <= 32'b000000_00110_00111_10110_00000_000010; 	// mul
		disk[1777] <= 32'b010010_11110_10110_1111111111111111; 	// sw
		disk[1778] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1779] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[1780] <= 32'b000000_00101_01111_10111_00000_010000; 	// gt
		disk[1781] <= 32'b010101_10111_00000_0000011100001001; 	// jf
		disk[1782] <= 32'b001111_11110_00110_1111111111111110; 	// lw
		disk[1783] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[1784] <= 32'b001111_00001_10000_0000000000000000; 	// lw
		disk[1785] <= 32'b010010_11110_10000_1111111111111101; 	// sw
		disk[1786] <= 32'b001111_11110_00111_1111111111111101; 	// lw
		disk[1787] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[1788] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[1789] <= 32'b001110_01000_00010_0000000000000000; 	// mov
		disk[1790] <= 32'b010010_00010_00001_0000000000000000; 	// sw
		disk[1791] <= 32'b000001_00110_10001_0000000000000001; 	// addi
		disk[1792] <= 32'b010010_11110_10001_1111111111111110; 	// sw
		disk[1793] <= 32'b001111_11110_00110_1111111111111110; 	// lw
		disk[1794] <= 32'b000001_01000_10010_0000000000000001; 	// addi
		disk[1795] <= 32'b010010_11110_10010_1111111111111111; 	// sw
		disk[1796] <= 32'b001111_11110_01000_1111111111111111; 	// lw
		disk[1797] <= 32'b000010_00101_10011_0000000000000001; 	// subi
		disk[1798] <= 32'b010010_11110_10011_0000000000000000; 	// sw
		disk[1799] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1800] <= 32'b111100_00000000000000011011110010; 	// j
		disk[1801] <= 32'b001111_11110_00101_1111111111111100; 	// lw
		disk[1802] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1803] <= 32'b111110_00000000000000000001100011; 	// jal
		disk[1804] <= 32'b000010_11110_11110_0000000000000110; 	// subi
		disk[1805] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1806] <= 32'b010001_11101_00110_0000000000000100; 	// la
		disk[1807] <= 32'b001111_11101_00111_0000000001011111; 	// lw
		disk[1808] <= 32'b000000_00110_00111_10100_00000_000000; 	// add
		disk[1809] <= 32'b001111_11101_01000_0000000000000001; 	// lw
		disk[1810] <= 32'b010010_10100_01000_0000000000000000; 	// sw
		disk[1811] <= 32'b001111_11101_01001_0000000110101011; 	// lw
		disk[1812] <= 32'b010010_11101_01001_0000000110111101; 	// sw
		disk[1813] <= 32'b001111_11101_01010_0000000110111101; 	// lw
		disk[1814] <= 32'b001110_01010_00001_0000000000000000; 	// mov
		disk[1815] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[1816] <= 32'b010000_00000_11101_0000000000000000; 	// li
		disk[1817] <= 32'b010000_00000_11110_0000000111000111; 	// li
		disk[1818] <= 32'b100110_00000_00000_0000000000000000; 	// cic
		disk[1819] <= 32'b000001_00111_10101_0000000000000001; 	// addi
		disk[1820] <= 32'b001110_10101_00001_0000000000000000; 	// mov
		disk[1821] <= 32'b111110_00000000000000001111011001; 	// jal
		disk[1822] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[1823] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1824] <= 32'b111110_00000000000000010111011111; 	// jal
		disk[1825] <= 32'b000010_11110_11110_0000000000000011; 	// subi
		disk[1826] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1827] <= 32'b001111_11101_00110_0000000110101011; 	// lw
		disk[1828] <= 32'b010010_11101_00110_0000000110111101; 	// sw
		disk[1829] <= 32'b001111_11101_00111_0000000110111101; 	// lw
		disk[1830] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[1831] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[1832] <= 32'b010000_00000_11101_0000000000000000; 	// li
		disk[1833] <= 32'b010000_00000_11110_0000000111000111; 	// li
		disk[1834] <= 32'b100110_00000_00000_0000000000000000; 	// cic
		disk[1835] <= 32'b010000_00000_10110_0000000000000001; 	// li
		disk[1836] <= 32'b010101_10110_00000_0000100000110000; 	// jf
		disk[1837] <= 32'b010011_00000_10111_0000000000000000; 	// in
		disk[1838] <= 32'b010010_11110_10111_1111111111111001; 	// sw
		disk[1839] <= 32'b001111_11101_00101_0000000110111101; 	// lw
		disk[1840] <= 32'b001111_11101_00110_0000000110101011; 	// lw
		disk[1841] <= 32'b000000_00101_00110_01111_00000_001100; 	// eq
		disk[1842] <= 32'b010101_01111_00000_0000011101011000; 	// jf
		disk[1843] <= 32'b001111_11110_00111_1111111111111001; 	// lw
		disk[1844] <= 32'b010000_00000_10001_0000000000000001; 	// li
		disk[1845] <= 32'b000000_00111_10001_10000_00000_001100; 	// eq
		disk[1846] <= 32'b010101_10000_00000_0000011100111011; 	// jf
		disk[1847] <= 32'b001111_11101_01000_0000000110101100; 	// lw
		disk[1848] <= 32'b010010_11110_01000_1111111111111001; 	// sw
		disk[1849] <= 32'b001111_11110_00111_1111111111111001; 	// lw
		disk[1850] <= 32'b111100_00000000000000011101010111; 	// j
		disk[1851] <= 32'b001111_11110_00101_1111111111111001; 	// lw
		disk[1852] <= 32'b010000_00000_10011_0000000000000010; 	// li
		disk[1853] <= 32'b000000_00101_10011_10010_00000_001100; 	// eq
		disk[1854] <= 32'b010101_10010_00000_0000011101000011; 	// jf
		disk[1855] <= 32'b001111_11101_00110_0000000110110110; 	// lw
		disk[1856] <= 32'b010010_11110_00110_1111111111111001; 	// sw
		disk[1857] <= 32'b001111_11110_00101_1111111111111001; 	// lw
		disk[1858] <= 32'b111100_00000000000000011101010111; 	// j
		disk[1859] <= 32'b001111_11110_00101_1111111111111001; 	// lw
		disk[1860] <= 32'b010000_00000_10101_0000000000000011; 	// li
		disk[1861] <= 32'b000000_00101_10101_10100_00000_001100; 	// eq
		disk[1862] <= 32'b010101_10100_00000_0000011101001011; 	// jf
		disk[1863] <= 32'b001111_11101_00110_0000000110111001; 	// lw
		disk[1864] <= 32'b010010_11110_00110_1111111111111001; 	// sw
		disk[1865] <= 32'b001111_11110_00101_1111111111111001; 	// lw
		disk[1866] <= 32'b111100_00000000000000011101010111; 	// j
		disk[1867] <= 32'b001111_11110_00101_1111111111111001; 	// lw
		disk[1868] <= 32'b010000_00000_10111_0000000000000100; 	// li
		disk[1869] <= 32'b000000_00101_10111_10110_00000_001100; 	// eq
		disk[1870] <= 32'b010101_10110_00000_0000011101010101; 	// jf
		disk[1871] <= 32'b111110_00000000000000000000110011; 	// jal
		disk[1872] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[1873] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1874] <= 32'b001111_11101_00110_0000000110101011; 	// lw
		disk[1875] <= 32'b010010_11110_00110_1111111111111001; 	// sw
		disk[1876] <= 32'b111100_00000000000000011101010111; 	// j
		disk[1877] <= 32'b001111_11101_00101_0000000110101011; 	// lw
		disk[1878] <= 32'b010010_11110_00101_1111111111111001; 	// sw
		disk[1879] <= 32'b111100_00000000000000100000101010; 	// j
		disk[1880] <= 32'b001111_11101_00101_0000000110111101; 	// lw
		disk[1881] <= 32'b001111_11101_00110_0000000110101100; 	// lw
		disk[1882] <= 32'b000000_00101_00110_01111_00000_001100; 	// eq
		disk[1883] <= 32'b010101_01111_00000_0000011110000011; 	// jf
		disk[1884] <= 32'b001111_11110_00111_1111111111111001; 	// lw
		disk[1885] <= 32'b010000_00000_10001_0000000000000001; 	// li
		disk[1886] <= 32'b000000_00111_10001_10000_00000_001100; 	// eq
		disk[1887] <= 32'b010101_10000_00000_0000011101100110; 	// jf
		disk[1888] <= 32'b111110_00000000000000010010001101; 	// jal
		disk[1889] <= 32'b000010_11110_11110_0000000000000110; 	// subi
		disk[1890] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1891] <= 32'b001111_11101_00110_0000000110101011; 	// lw
		disk[1892] <= 32'b010010_11110_00110_1111111111111001; 	// sw
		disk[1893] <= 32'b111100_00000000000000011110000010; 	// j
		disk[1894] <= 32'b001111_11110_00101_1111111111111001; 	// lw
		disk[1895] <= 32'b010000_00000_10011_0000000000000010; 	// li
		disk[1896] <= 32'b000000_00101_10011_10010_00000_001100; 	// eq
		disk[1897] <= 32'b010101_10010_00000_0000011101110011; 	// jf
		disk[1898] <= 32'b001111_11101_00110_0000000110101110; 	// lw
		disk[1899] <= 32'b010010_11110_00110_1111111111111001; 	// sw
		disk[1900] <= 32'b001111_11110_00101_1111111111111001; 	// lw
		disk[1901] <= 32'b111110_00000000000000000100111101; 	// jal
		disk[1902] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[1903] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1904] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1905] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
		disk[1906] <= 32'b111100_00000000000000011110000010; 	// j
		disk[1907] <= 32'b001111_11110_00101_1111111111111001; 	// lw
		disk[1908] <= 32'b010000_00000_10101_0000000000000011; 	// li
		disk[1909] <= 32'b000000_00101_10101_10100_00000_001100; 	// eq
		disk[1910] <= 32'b010101_10100_00000_0000011110000000; 	// jf
		disk[1911] <= 32'b001111_11101_00110_0000000110101101; 	// lw
		disk[1912] <= 32'b010010_11110_00110_1111111111111001; 	// sw
		disk[1913] <= 32'b001111_11110_00101_1111111111111001; 	// lw
		disk[1914] <= 32'b111110_00000000000000000100111101; 	// jal
		disk[1915] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[1916] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1917] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1918] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
		disk[1919] <= 32'b111100_00000000000000011110000010; 	// j
		disk[1920] <= 32'b001111_11101_00101_0000000110101011; 	// lw
		disk[1921] <= 32'b010010_11110_00101_1111111111111001; 	// sw
		disk[1922] <= 32'b111100_00000000000000100000101010; 	// j
		disk[1923] <= 32'b001111_11101_00101_0000000110111101; 	// lw
		disk[1924] <= 32'b001111_11101_00110_0000000110101101; 	// lw
		disk[1925] <= 32'b000000_00101_00110_10110_00000_001100; 	// eq
		disk[1926] <= 32'b010101_10110_00000_0000011110010010; 	// jf
		disk[1927] <= 32'b001111_11110_00111_1111111111111001; 	// lw
		disk[1928] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[1929] <= 32'b000000_00111_01111_10111_00000_010000; 	// gt
		disk[1930] <= 32'b010101_10111_00000_0000011110001111; 	// jf
		disk[1931] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[1932] <= 32'b111110_00000000000000000011101001; 	// jal
		disk[1933] <= 32'b000010_11110_11110_0000000000000101; 	// subi
		disk[1934] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1935] <= 32'b001111_11101_00101_0000000110101011; 	// lw
		disk[1936] <= 32'b010010_11110_00101_1111111111111001; 	// sw
		disk[1937] <= 32'b111100_00000000000000100000101010; 	// j
		disk[1938] <= 32'b001111_11101_00101_0000000110111101; 	// lw
		disk[1939] <= 32'b001111_11101_00110_0000000110101110; 	// lw
		disk[1940] <= 32'b000000_00101_00110_10000_00000_001100; 	// eq
		disk[1941] <= 32'b010101_10000_00000_0000011110100001; 	// jf
		disk[1942] <= 32'b001111_11110_00111_1111111111111001; 	// lw
		disk[1943] <= 32'b010000_00000_10010_0000000000000000; 	// li
		disk[1944] <= 32'b000000_00111_10010_10001_00000_010000; 	// gt
		disk[1945] <= 32'b010101_10001_00000_0000011110011110; 	// jf
		disk[1946] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[1947] <= 32'b111110_00000000000000000100101101; 	// jal
		disk[1948] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[1949] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1950] <= 32'b001111_11101_00101_0000000110101011; 	// lw
		disk[1951] <= 32'b010010_11110_00101_1111111111111001; 	// sw
		disk[1952] <= 32'b111100_00000000000000100000101010; 	// j
		disk[1953] <= 32'b001111_11101_00101_0000000110111101; 	// lw
		disk[1954] <= 32'b001111_11101_00110_0000000110110110; 	// lw
		disk[1955] <= 32'b000000_00101_00110_10011_00000_001100; 	// eq
		disk[1956] <= 32'b010101_10011_00000_0000011111000010; 	// jf
		disk[1957] <= 32'b001111_11110_00111_1111111111111001; 	// lw
		disk[1958] <= 32'b010000_00000_10101_0000000000000001; 	// li
		disk[1959] <= 32'b000000_00111_10101_10100_00000_001100; 	// eq
		disk[1960] <= 32'b010101_10100_00000_0000011110110010; 	// jf
		disk[1961] <= 32'b001111_11101_01000_0000000110110111; 	// lw
		disk[1962] <= 32'b010010_11110_01000_1111111111111001; 	// sw
		disk[1963] <= 32'b001111_11110_00111_1111111111111001; 	// lw
		disk[1964] <= 32'b111110_00000000000000000100111101; 	// jal
		disk[1965] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[1966] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1967] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1968] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
		disk[1969] <= 32'b111100_00000000000000011111000001; 	// j
		disk[1970] <= 32'b001111_11110_00101_1111111111111001; 	// lw
		disk[1971] <= 32'b010000_00000_10111_0000000000000010; 	// li
		disk[1972] <= 32'b000000_00101_10111_10110_00000_001100; 	// eq
		disk[1973] <= 32'b010101_10110_00000_0000011110111111; 	// jf
		disk[1974] <= 32'b001111_11101_00110_0000000110111000; 	// lw
		disk[1975] <= 32'b010010_11110_00110_1111111111111001; 	// sw
		disk[1976] <= 32'b001111_11110_00101_1111111111111001; 	// lw
		disk[1977] <= 32'b111110_00000000000000000101100010; 	// jal
		disk[1978] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[1979] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1980] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1981] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
		disk[1982] <= 32'b111100_00000000000000011111000001; 	// j
		disk[1983] <= 32'b001111_11101_00101_0000000110101011; 	// lw
		disk[1984] <= 32'b010010_11110_00101_1111111111111001; 	// sw
		disk[1985] <= 32'b111100_00000000000000100000101010; 	// j
		disk[1986] <= 32'b001111_11101_00101_0000000110111101; 	// lw
		disk[1987] <= 32'b001111_11101_00110_0000000110110111; 	// lw
		disk[1988] <= 32'b000000_00101_00110_01111_00000_001100; 	// eq
		disk[1989] <= 32'b010101_01111_00000_0000011111010001; 	// jf
		disk[1990] <= 32'b001111_11110_00111_1111111111111001; 	// lw
		disk[1991] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[1992] <= 32'b000000_00111_10001_10000_00000_010000; 	// gt
		disk[1993] <= 32'b010101_10000_00000_0000011111001110; 	// jf
		disk[1994] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[1995] <= 32'b111110_00000000000000010000101111; 	// jal
		disk[1996] <= 32'b000010_11110_11110_0000000000001010; 	// subi
		disk[1997] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[1998] <= 32'b001111_11101_00101_0000000110101011; 	// lw
		disk[1999] <= 32'b010010_11110_00101_1111111111111001; 	// sw
		disk[2000] <= 32'b111100_00000000000000100000101010; 	// j
		disk[2001] <= 32'b001111_11101_00101_0000000110111101; 	// lw
		disk[2002] <= 32'b001111_11101_00110_0000000110111000; 	// lw
		disk[2003] <= 32'b000000_00101_00110_10010_00000_001100; 	// eq
		disk[2004] <= 32'b010101_10010_00000_0000011111100000; 	// jf
		disk[2005] <= 32'b001111_11110_00111_1111111111111001; 	// lw
		disk[2006] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[2007] <= 32'b000000_00111_10100_10011_00000_010000; 	// gt
		disk[2008] <= 32'b010101_10011_00000_0000011111011101; 	// jf
		disk[2009] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[2010] <= 32'b111110_00000000000000000010100000; 	// jal
		disk[2011] <= 32'b000010_11110_11110_0000000000000101; 	// subi
		disk[2012] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[2013] <= 32'b001111_11101_00101_0000000110101011; 	// lw
		disk[2014] <= 32'b010010_11110_00101_1111111111111001; 	// sw
		disk[2015] <= 32'b111100_00000000000000100000101010; 	// j
		disk[2016] <= 32'b001111_11101_00101_0000000110111101; 	// lw
		disk[2017] <= 32'b001111_11101_00110_0000000110111001; 	// lw
		disk[2018] <= 32'b000000_00101_00110_10101_00000_001100; 	// eq
		disk[2019] <= 32'b010101_10101_00000_0000100000001011; 	// jf
		disk[2020] <= 32'b001111_11110_00111_1111111111111001; 	// lw
		disk[2021] <= 32'b010000_00000_10111_0000000000000001; 	// li
		disk[2022] <= 32'b000000_00111_10111_10110_00000_001100; 	// eq
		disk[2023] <= 32'b010101_10110_00000_0000011111110000; 	// jf
		disk[2024] <= 32'b010000_00000_01111_0000000000000001; 	// li
		disk[2025] <= 32'b010010_11101_01111_0000000001101010; 	// sw
		disk[2026] <= 32'b111110_00000000000000010111011111; 	// jal
		disk[2027] <= 32'b000010_11110_11110_0000000000000011; 	// subi
		disk[2028] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[2029] <= 32'b001111_11101_00110_0000000110101011; 	// lw
		disk[2030] <= 32'b010010_11110_00110_1111111111111001; 	// sw
		disk[2031] <= 32'b111100_00000000000000100000001010; 	// j
		disk[2032] <= 32'b001111_11110_00101_1111111111111001; 	// lw
		disk[2033] <= 32'b010000_00000_10001_0000000000000010; 	// li
		disk[2034] <= 32'b000000_00101_10001_10000_00000_001100; 	// eq
		disk[2035] <= 32'b010101_10000_00000_0000011111111100; 	// jf
		disk[2036] <= 32'b111110_00000000000000000101100010; 	// jal
		disk[2037] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[2038] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[2039] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[2040] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
		disk[2041] <= 32'b001111_11101_00110_0000000110111010; 	// lw
		disk[2042] <= 32'b010010_11110_00110_1111111111111001; 	// sw
		disk[2043] <= 32'b111100_00000000000000100000001010; 	// j
		disk[2044] <= 32'b001111_11110_00101_1111111111111001; 	// lw
		disk[2045] <= 32'b010000_00000_10011_0000000000000011; 	// li
		disk[2046] <= 32'b000000_00101_10011_10010_00000_001100; 	// eq
		disk[2047] <= 32'b010101_10010_00000_0000100000001000; 	// jf
		disk[2048] <= 32'b111110_00000000000000000110000111; 	// jal
		disk[2049] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[2050] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[2051] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[2052] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
		disk[2053] <= 32'b001111_11101_00110_0000000110111011; 	// lw
		disk[2054] <= 32'b010010_11110_00110_1111111111111001; 	// sw
		disk[2055] <= 32'b111100_00000000000000100000001010; 	// j
		disk[2056] <= 32'b001111_11101_00101_0000000110101011; 	// lw
		disk[2057] <= 32'b010010_11110_00101_1111111111111001; 	// sw
		disk[2058] <= 32'b111100_00000000000000100000101010; 	// j
		disk[2059] <= 32'b001111_11101_00101_0000000110111101; 	// lw
		disk[2060] <= 32'b001111_11101_00110_0000000110111010; 	// lw
		disk[2061] <= 32'b000000_00101_00110_10100_00000_001100; 	// eq
		disk[2062] <= 32'b010101_10100_00000_0000100000011100; 	// jf
		disk[2063] <= 32'b001111_11110_00111_1111111111111001; 	// lw
		disk[2064] <= 32'b010000_00000_10110_0000000000000000; 	// li
		disk[2065] <= 32'b000000_00111_10110_10101_00000_010000; 	// gt
		disk[2066] <= 32'b010101_10101_00000_0000100000011001; 	// jf
		disk[2067] <= 32'b010000_00000_10111_0000000000000000; 	// li
		disk[2068] <= 32'b010010_11101_10111_0000000001101010; 	// sw
		disk[2069] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[2070] <= 32'b111110_00000000000000010111001001; 	// jal
		disk[2071] <= 32'b000010_11110_11110_0000000000000011; 	// subi
		disk[2072] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[2073] <= 32'b001111_11101_00101_0000000110101011; 	// lw
		disk[2074] <= 32'b010010_11110_00101_1111111111111001; 	// sw
		disk[2075] <= 32'b111100_00000000000000100000101010; 	// j
		disk[2076] <= 32'b001111_11101_00101_0000000110111101; 	// lw
		disk[2077] <= 32'b001111_11101_00110_0000000110111011; 	// lw
		disk[2078] <= 32'b000000_00101_00110_01111_00000_001100; 	// eq
		disk[2079] <= 32'b010101_01111_00000_0000100000101010; 	// jf
		disk[2080] <= 32'b001111_11110_00111_1111111111111001; 	// lw
		disk[2081] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[2082] <= 32'b000000_00111_10001_10000_00000_010000; 	// gt
		disk[2083] <= 32'b010101_10000_00000_0000100000101000; 	// jf
		disk[2084] <= 32'b001110_00111_00001_0000000000000000; 	// mov
		disk[2085] <= 32'b111110_00000000000000010110101110; 	// jal
		disk[2086] <= 32'b000010_11110_11110_0000000000000011; 	// subi
		disk[2087] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[2088] <= 32'b001111_11101_00101_0000000110101011; 	// lw
		disk[2089] <= 32'b010010_11110_00101_1111111111111001; 	// sw
		disk[2090] <= 32'b001111_11110_00101_1111111111111001; 	// lw
		disk[2091] <= 32'b010010_11101_00101_0000000110111101; 	// sw
		disk[2092] <= 32'b001111_11101_00110_0000000110111101; 	// lw
		disk[2093] <= 32'b001110_00110_00001_0000000000000000; 	// mov
		disk[2094] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
		disk[2095] <= 32'b111100_00000000000000011100101011; 	// j
		disk[2096] <= 32'b111111_00000000000000000000000000; 	// halt

		// PROGRAMA 1
		disk[3800] <= 32'b111101_00000000000000000000100011;		// Jump to Main
		disk[3801] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[3802] <= 32'b010010_11110_00001_1111111111111100; 	// sw
		disk[3803] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[3804] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[3805] <= 32'b010000_00000_10000_0000000000000001; 	// li
		disk[3806] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[3807] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[3808] <= 32'b010010_11110_10001_1111111111111101; 	// sw
		disk[3809] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[3810] <= 32'b001111_11110_00110_1111111111111100; 	// lw
		disk[3811] <= 32'b000000_00101_00110_10010_00000_001111; 	// let
		disk[3812] <= 32'b010101_10010_00000_0000000000100000; 	// jf
		disk[3813] <= 32'b010000_00000_10100_0000000000000001; 	// li
		disk[3814] <= 32'b000000_00101_10100_10011_00000_001111; 	// let
		disk[3815] <= 32'b010101_10011_00000_0000000000010010; 	// jf
		disk[3816] <= 32'b010010_11110_00101_1111111111111110; 	// sw
		disk[3817] <= 32'b111100_00000000000000000000011011; 	// j
		disk[3818] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[3819] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[3820] <= 32'b000000_00101_00110_10101_00000_000000; 	// add
		disk[3821] <= 32'b010010_11110_10101_1111111111111110; 	// sw
		disk[3822] <= 32'b010010_11110_00110_1111111111111111; 	// sw
		disk[3823] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[3824] <= 32'b001111_11110_00111_1111111111111110; 	// lw
		disk[3825] <= 32'b010010_11110_00111_0000000000000000; 	// sw
		disk[3826] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[3827] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[3828] <= 32'b000001_00101_10110_0000000000000001; 	// addi
		disk[3829] <= 32'b010010_11110_10110_1111111111111101; 	// sw
		disk[3830] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[3831] <= 32'b111100_00000000000000000000001001; 	// j
		disk[3832] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[3833] <= 32'b001110_00101_11000_0000000000000000; 	// mov
		disk[3834] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[3835] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[3836] <= 32'b010000_00000_01111_0000000000001011; 	// li
		disk[3837] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[3838] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[3839] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[3840] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[3841] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[3842] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[3843] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[3844] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[3845] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[3846] <= 32'b010000_00000_00010_0000000000000000; 	// li
		disk[3847] <= 32'b010100_00000_00001_0000000000000000; 	// out
		disk[3848] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[3849] <= 32'b011111_11001_00000_0000000000000000; 	// syscall

		// PROGRAMA 2
		disk[3900] <= 32'b111101_00000000000000000000100001;		// Jump to Main
		disk[3901] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[3902] <= 32'b010010_11110_00001_1111111111111100; 	// sw
		disk[3903] <= 32'b010010_11110_00010_1111111111111101; 	// sw
		disk[3904] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[3905] <= 32'b010010_11110_01111_1111111111111110; 	// sw
		disk[3906] <= 32'b010000_00000_10000_0000000000000000; 	// li
		disk[3907] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[3908] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[3909] <= 32'b001111_11110_00110_1111111111111101; 	// lw
		disk[3910] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
		disk[3911] <= 32'b010101_10001_00000_0000000000011100; 	// jf
		disk[3912] <= 32'b001111_11110_00111_1111111111111100; 	// lw
		disk[3913] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
		disk[3914] <= 32'b001111_10010_10010_0000000000000000; 	// lw
		disk[3915] <= 32'b001111_11110_01000_0000000000000000; 	// lw
		disk[3916] <= 32'b000000_01000_10010_10011_00000_001110; 	// lt
		disk[3917] <= 32'b010101_10011_00000_0000000000010111; 	// jf
		disk[3918] <= 32'b000000_00111_00101_10100_00000_000000; 	// add
		disk[3919] <= 32'b001111_10100_10100_0000000000000000; 	// lw
		disk[3920] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[3921] <= 32'b001111_11110_01000_0000000000000000; 	// lw
		disk[3922] <= 32'b010010_11110_00101_1111111111111111; 	// sw
		disk[3923] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[3924] <= 32'b000001_00101_10101_0000000000000001; 	// addi
		disk[3925] <= 32'b010010_11110_10101_1111111111111110; 	// sw
		disk[3926] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[3927] <= 32'b111100_00000000000000000000001000; 	// j
		disk[3928] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[3929] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[3930] <= 32'b010000_00000_00010_0000000000000001; 	// li
		disk[3931] <= 32'b010100_00000_00001_0000000000000001; 	// out
		disk[3932] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[3933] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[3934] <= 32'b010001_11110_00101_1111111111111011; 	// la
		disk[3935] <= 32'b010000_00000_01111_0000000000001100; 	// li
		disk[3936] <= 32'b010010_00101_01111_0000000000000000; 	// sw
		disk[3937] <= 32'b010000_00000_10000_0000000000101001; 	// li
		disk[3938] <= 32'b010010_00101_10000_0000000000000001; 	// sw
		disk[3939] <= 32'b010000_00000_10001_0000000000010111; 	// li
		disk[3940] <= 32'b010010_00101_10001_0000000000000010; 	// sw
		disk[3941] <= 32'b010000_00000_10010_0000000001100010; 	// li
		disk[3942] <= 32'b010010_00101_10010_0000000000000011; 	// sw
		disk[3943] <= 32'b010000_00000_10011_0000000000100001; 	// li
		disk[3944] <= 32'b010010_00101_10011_0000000000000100; 	// sw
		disk[3945] <= 32'b010000_00000_10100_0000000000010101; 	// li
		disk[3946] <= 32'b010010_00101_10100_0000000000000101; 	// sw
		disk[3947] <= 32'b010001_11110_00001_1111111111111011; 	// la
		disk[3948] <= 32'b010000_00000_00010_0000000000000110; 	// li
		disk[3949] <= 32'b010010_11110_11111_1111111111111010; 	// sw
		disk[3950] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[3951] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[3952] <= 32'b001111_11110_11111_1111111111111010; 	// lw
		disk[3953] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[3954] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[3955] <= 32'b011111_11001_00000_0000000000000000; 	// syscall
		
		// PROGRAMA 3
		disk[4000] <= 32'b111101_00000000000000000000010100;		// Jump to Main
		disk[4001] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[4002] <= 32'b010010_11110_00001_1111111111111111; 	// sw
		disk[4003] <= 32'b010000_00000_01111_0000000000000001; 	// li
		disk[4004] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[4005] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[4006] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[4007] <= 32'b000000_00101_10001_10000_00000_010000; 	// gt
		disk[4008] <= 32'b010101_10000_00000_0000000000010001; 	// jf
		disk[4009] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[4010] <= 32'b000000_00110_00101_10010_00000_000010; 	// mul
		disk[4011] <= 32'b010010_11110_10010_0000000000000000; 	// sw
		disk[4012] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[4013] <= 32'b000010_00101_10011_0000000000000001; 	// subi
		disk[4014] <= 32'b010010_11110_10011_1111111111111111; 	// sw
		disk[4015] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[4016] <= 32'b111100_00000000000000000000000101; 	// j
		disk[4017] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[4018] <= 32'b001110_00101_11000_0000000000000000; 	// mov
		disk[4019] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[4020] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[4021] <= 32'b101000_00000000000000000000000000; 	// preIO
		disk[4022] <= 32'b010011_00000_01111_0000000000000000; 	// in
		disk[4023] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[4024] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[4025] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[4026] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[4027] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[4028] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[4029] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[4030] <= 32'b001110_11000_00101_0000000000000000; 	// mov
		disk[4031] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[4032] <= 32'b010000_00000_00010_0000000000000010; 	// li
		disk[4033] <= 32'b010100_00000_00001_0000000000000010; 	// out
		disk[4034] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[4035] <= 32'b011111_11001_00000_0000000000000000; 	// syscall
		
	end
endmodule
