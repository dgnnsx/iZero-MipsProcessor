library verilog;
use verilog.vl_types.all;
entity entrada_de_dados_vlg_vec_tst is
end entrada_de_dados_vlg_vec_tst;
