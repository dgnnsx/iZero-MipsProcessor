module disco_rigido (clk, we, addr, datain, dataout);
	input clk;										// clock
	input we;										// write enable
	input [31:0] addr;							// disk address
	input [31:0] datain;							// data in (to disk)
	
	output reg [31:0] dataout;					// data out (from disk)
	
	localparam DISK_SIZE = 100;				// Tamanho do disco
	reg [31:0] disk [DISK_SIZE-1:0];			// disk cells
	
	always @ (posedge clk) begin
		if (we) disk[addr] <= datain;			// write disk
	end
	
	always @ (negedge clk) begin
		dataout <= disk[addr];
	end

	initial begin
		disk[0] <= 32'b010110_00000000000000000000101110;		// Jump to Main
		disk[1] <= 32'b000001_11110_11110_0000000000001000; 	// addi
		disk[2] <= 32'b010010_11110_00110_1111111111111011; 	// sw
		disk[3] <= 32'b010010_11110_00111_1111111111111100; 	// sw
		disk[4] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[5] <= 32'b010010_11110_10100_1111111111111101; 	// sw
		disk[6] <= 32'b001111_11110_01010_1111111111111100; 	// lw
		disk[7] <= 32'b000010_01010_10101_0000000000000001; 	// subi
		disk[8] <= 32'b001111_11110_01011_1111111111111101; 	// lw
		disk[9] <= 32'b000000_01011_10101_10110_00000_001110; 	// lt
		disk[10] <= 32'b010101_10110_00000_0000000000101101; 	// jf
		disk[11] <= 32'b010010_11110_01011_1111111111111111; 	// sw
		disk[12] <= 32'b000001_01011_10111_0000000000000001; 	// addi
		disk[13] <= 32'b010010_11110_10111_1111111111111110; 	// sw
		disk[14] <= 32'b001111_11110_01100_1111111111111110; 	// lw
		disk[15] <= 32'b000000_01100_01010_11000_00000_001110; 	// lt
		disk[16] <= 32'b010101_11000_00000_0000000000011101; 	// jf
		disk[17] <= 32'b001111_11110_01101_1111111111111011; 	// lw
		disk[18] <= 32'b000000_01101_01100_11001_00000_000000; 	// add
		disk[19] <= 32'b001111_11001_11001_0000000000000000; 	// lw
		disk[20] <= 32'b001111_11110_01110_1111111111111111; 	// lw
		disk[21] <= 32'b000000_01101_01110_11010_00000_000000; 	// add
		disk[22] <= 32'b001111_11010_11010_0000000000000000; 	// lw
		disk[23] <= 32'b000000_11001_11010_11011_00000_001110; 	// lt
		disk[24] <= 32'b010101_11011_00000_0000000000011010; 	// jf
		disk[25] <= 32'b010010_11110_01100_1111111111111111; 	// sw
		disk[26] <= 32'b000001_01100_11100_0000000000000001; 	// addi
		disk[27] <= 32'b010010_11110_11100_1111111111111110; 	// sw
		disk[28] <= 32'b010110_00000000000000000000001110; 	// j
		disk[29] <= 32'b001111_11110_01111_1111111111111111; 	// lw
		disk[30] <= 32'b000000_01011_01111_11101_00000_001101; 	// ne
		disk[31] <= 32'b010101_11101_00000_0000000000101010; 	// jf
		disk[32] <= 32'b000000_01101_01011_10100_00000_000000; 	// add
		disk[33] <= 32'b001111_10100_10100_0000000000000000; 	// lw
		disk[34] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[35] <= 32'b000000_01101_01111_10101_00000_000000; 	// add
		disk[36] <= 32'b001111_10101_10101_0000000000000000; 	// lw
		disk[37] <= 32'b000000_01101_01011_10110_00000_000000; 	// add
		disk[38] <= 32'b010010_10110_10101_0000000000000000; 	// sw
		disk[39] <= 32'b000000_01101_01111_10111_00000_000000; 	// add
		disk[40] <= 32'b001111_11110_10000_0000000000000000; 	// lw
		disk[41] <= 32'b010010_10111_10000_0000000000000000; 	// sw
		disk[42] <= 32'b000001_01011_11000_0000000000000001; 	// addi
		disk[43] <= 32'b010010_11110_11000_1111111111111101; 	// sw
		disk[44] <= 32'b010110_00000000000000000000000110; 	// j
		disk[45] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[46] <= 32'b000001_11110_11110_0000000000000101; 	// addi
		disk[47] <= 32'b010001_11110_01010_1111111111111100; 	// la
		disk[48] <= 32'b010000_00000_10100_0000000000001001; 	// li
		disk[49] <= 32'b010010_01010_10100_0000000000000000; 	// sw
		disk[50] <= 32'b010000_00000_10101_0000000000000110; 	// li
		disk[51] <= 32'b010010_01010_10101_0000000000000001; 	// sw
		disk[52] <= 32'b010000_00000_10110_0000000000001000; 	// li
		disk[53] <= 32'b010010_01010_10110_0000000000000010; 	// sw
		disk[54] <= 32'b010000_00000_10111_0000000000000111; 	// li
		disk[55] <= 32'b010010_01010_10111_0000000000000011; 	// sw
		disk[56] <= 32'b010001_11110_00110_1111111111111100; 	// la
		disk[57] <= 32'b010000_00000_00111_0000000000000100; 	// li
		disk[58] <= 32'b010111_00000000000000000000000001; 	// jal
		disk[59] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[60] <= 32'b000010_11110_11110_0000000000001000; 	// subi
		disk[61] <= 32'b010011_00000_11000_0000000000000000; 	// in
		disk[62] <= 32'b010010_11110_11000_0000000000000000; 	// sw
		disk[63] <= 32'b010001_11110_01100_1111111111111100; 	// la
		disk[64] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[65] <= 32'b000000_01100_01101_11001_00000_000000; 	// add
		disk[66] <= 32'b001111_11001_11001_0000000000000000; 	// lw
		disk[67] <= 32'b001110_11001_00110_0000000000000000; 	// mov
		disk[68] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[69] <= 32'b010100_00000_00110_0000000000000010; 	// out
		disk[70] <= 32'b011000_00000000000000000000000000; 	// halt
	end
endmodule
