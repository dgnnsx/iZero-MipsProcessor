library verilog;
use verilog.vl_types.all;
entity saida_de_dados_vlg_vec_tst is
end saida_de_dados_vlg_vec_tst;
