library verilog;
use verilog.vl_types.all;
entity extensor_de_bit_vlg_vec_tst is
end extensor_de_bit_vlg_vec_tst;
