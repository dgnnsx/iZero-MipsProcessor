module memoria_de_instrucoes(pc, instrucao);
	// Entrada
	input [25:0] pc;				// PC Atual
	
	// Saida
	output [31:0] instrucao;	// Proxima instrucao a ser executada
	
	parameter MEM_SIZE = 150; // Tamanho da memoria
	wire [31:0] rom [MEM_SIZE-1:0];// Memoria de instrucoes

assign rom[0] = 32'b010110_00000000000000000000011110;		// Jump to Main
assign rom[1] = 32'b000001_00011_00011_0000000000000110; 	// addi
assign rom[2] = 32'b010010_00011_00111_1111111111111100; 	// sw
assign rom[3] = 32'b010000_00000_10101_0000000000000000; 	// li
assign rom[4] = 32'b010010_00011_10101_1111111111111111; 	// sw
assign rom[5] = 32'b010000_00000_10110_0000000000000001; 	// li
assign rom[6] = 32'b010010_00011_10110_0000000000000000; 	// sw
assign rom[7] = 32'b010000_00000_10111_0000000000000000; 	// li
assign rom[8] = 32'b010010_00011_10111_1111111111111101; 	// sw
assign rom[9] = 32'b001111_00011_01011_1111111111111101; 	// lw
assign rom[10] = 32'b001111_00011_01100_1111111111111100; 	// lw
assign rom[11] = 32'b000000_01011_01100_11000_00000_001111; 	// get
assign rom[12] = 32'b010101_11000_00000_0000000000011100; 	// jf
assign rom[13] = 32'b010000_00000_11010_0000000000000001; 	// li
assign rom[14] = 32'b000000_01011_11010_11001_00000_001111; 	// get
assign rom[15] = 32'b010101_11001_00000_0000000000010010; 	// jf
assign rom[16] = 32'b010010_00011_01011_1111111111111110; 	// sw
assign rom[17] = 32'b010110_00000000000000000000011001; 	// j
assign rom[18] = 32'b001111_00011_01101_1111111111111111; 	// lw
assign rom[19] = 32'b001111_00011_01110_0000000000000000; 	// lw
assign rom[20] = 32'b000000_01101_01110_11011_00000_000000; 	// add
assign rom[21] = 32'b010010_00011_11011_1111111111111110; 	// sw
assign rom[22] = 32'b010010_00011_01110_1111111111111111; 	// sw
assign rom[23] = 32'b001111_00011_01111_1111111111111110; 	// lw
assign rom[24] = 32'b010010_00011_01111_0000000000000000; 	// sw
assign rom[25] = 32'b000001_01011_11100_0000000000000001; 	// addi
assign rom[26] = 32'b010010_00011_11100_1111111111111101; 	// sw
assign rom[27] = 32'b010110_00000000000000000000001001; 	// j
assign rom[28] = 32'b001110_01111_00001_0000000000000000; 	// mov
assign rom[29] = 32'b000000_11111_00000_00000_00000_010010; 	// jr
assign rom[30] = 32'b000001_00011_00011_0000000000000001; 	// addi
assign rom[31] = 32'b010011_00000_10101_0000000000000000; 	// in
assign rom[32] = 32'b010010_00011_10101_0000000000000000; 	// sw
assign rom[33] = 32'b001111_00011_01011_0000000000000000; 	// lw
assign rom[34] = 32'b001110_01011_00111_0000000000000000; 	// mov
assign rom[35] = 32'b010111_00000000000000000000000001; 	// jal
assign rom[36] = 32'b001110_00001_10110_0000000000000000; 	// mov
assign rom[37] = 32'b000010_00011_00011_0000000000000110; 	// subi
assign rom[38] = 32'b001110_10110_00111_0000000000000000; 	// mov
assign rom[39] = 32'b010000_00000_01000_0000000000000010; 	// li
assign rom[40] = 32'b010100_00000_00111_0000000000000010; 	// out
assign rom[41] = 32'b011000_00000000000000000000000000; 	// halt
	
	assign instrucao = rom[pc];
endmodule
