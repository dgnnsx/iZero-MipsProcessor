module disco_rigido (clk, we, addr, datain, dataout);
	input clk;										// clock
	input we;										// write enable
	input [31:0] addr;							// disk address
	input [31:0] datain;							// data in (to disk)
	
	output reg [31:0] dataout;					// data out (from disk)
	
	localparam DISK_SIZE = 1024;				// Tamanho do disco
	reg [31:0] disk [DISK_SIZE-1:0];			// disk cells
	
	always @ (posedge clk) begin
		if (we) disk[addr] <= datain;			// write disk
	end
	
	always @ (negedge clk) begin
		dataout <= disk[addr];
	end

	initial begin
		// SISTEMA OPERACIONAL

		disk[0] <= 32'b010110_00000000000000000000000001;		// Jump to Main
disk[1] <= 32'b001110_00000_00101_0000000000000000; 	// mov
disk[2] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[3] <= 32'b010000_00000_10100_0000000000010100; 	// li
disk[4] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[5] <= 32'b010000_00000_10101_0000000000011110; 	// li
disk[6] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[7] <= 32'b001111_11110_01010_1111111111111111; 	// lw
disk[8] <= 32'b010000_00000_10111_0000000000001010; 	// li
disk[9] <= 32'b000000_01010_10111_10110_00000_010000; 	// gt
disk[10] <= 32'b001111_11110_01011_0000000000000000; 	// lw
disk[11] <= 32'b010000_00000_11001_0000000000001010; 	// li
disk[12] <= 32'b000000_01011_11001_11000_00000_010000; 	// gt
disk[13] <= 32'b000000_10110_11000_11010_00000_001000; 	// land
disk[14] <= 32'b010101_11010_00000_0000000000010011; 	// jf
disk[15] <= 32'b010000_00000_00110_0000000000001011; 	// li
disk[16] <= 32'b010000_00000_00111_0000000000000000; 	// li
disk[17] <= 32'b010100_00000_00110_0000000000000000; 	// out
disk[18] <= 32'b010110_00000000000000000000010110; 	// j
disk[19] <= 32'b010000_00000_00110_0000000000010110; 	// li
disk[20] <= 32'b010000_00000_00111_0000000000000000; 	// li
disk[21] <= 32'b010100_00000_00110_0000000000000000; 	// out
disk[22] <= 32'b010000_00000_11100_0000000000010100; 	// li
disk[23] <= 32'b000000_01010_11100_11011_00000_010000; 	// gt
disk[24] <= 32'b010000_00000_10100_0000000000010100; 	// li
disk[25] <= 32'b000000_01011_10100_11101_00000_010000; 	// gt
disk[26] <= 32'b000000_11011_11101_10101_00000_001000; 	// land
disk[27] <= 32'b010101_10101_00000_0000000000100000; 	// jf
disk[28] <= 32'b010000_00000_00110_0000000000001011; 	// li
disk[29] <= 32'b010000_00000_00111_0000000000000001; 	// li
disk[30] <= 32'b010100_00000_00110_0000000000000001; 	// out
disk[31] <= 32'b010110_00000000000000000000100011; 	// j
disk[32] <= 32'b010000_00000_00110_0000000000010110; 	// li
disk[33] <= 32'b010000_00000_00111_0000000000000001; 	// li
disk[34] <= 32'b010100_00000_00110_0000000000000001; 	// out
disk[35] <= 32'b011000_00000000000000000000000000; 	// halt

		
		// PROGRAMA 1
		disk[800] <= 32'b010110_00000000000000000000100001;		// Jump to Main
		disk[801] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[802] <= 32'b010010_11110_00110_1111111111111100; 	// sw
		disk[803] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[804] <= 32'b010010_11110_10100_1111111111111111; 	// sw
		disk[805] <= 32'b010000_00000_10101_0000000000000001; 	// li
		disk[806] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[807] <= 32'b010000_00000_10110_0000000000000000; 	// li
		disk[808] <= 32'b010010_11110_10110_1111111111111101; 	// sw
		disk[809] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[810] <= 32'b001111_11110_01011_1111111111111100; 	// lw
		disk[811] <= 32'b000000_01010_01011_10111_00000_001111; 	// let
		disk[812] <= 32'b010101_10111_00000_0000000000011111; 	// jf
		disk[813] <= 32'b010000_00000_11001_0000000000000001; 	// li
		disk[814] <= 32'b000000_01010_11001_11000_00000_001111; 	// let
		disk[815] <= 32'b010101_11000_00000_0000000000010010; 	// jf
		disk[816] <= 32'b010010_11110_01010_1111111111111110; 	// sw
		disk[817] <= 32'b010110_00000000000000000000011011; 	// j
		disk[818] <= 32'b001111_11110_01100_1111111111111111; 	// lw
		disk[819] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[820] <= 32'b000000_01100_01101_11010_00000_000000; 	// add
		disk[821] <= 32'b010010_11110_11010_1111111111111110; 	// sw
		disk[822] <= 32'b010010_11110_01101_1111111111111111; 	// sw
		disk[823] <= 32'b001111_11110_01100_1111111111111111; 	// lw
		disk[824] <= 32'b001111_11110_01110_1111111111111110; 	// lw
		disk[825] <= 32'b010010_11110_01110_0000000000000000; 	// sw
		disk[826] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[827] <= 32'b000001_01010_11011_0000000000000001; 	// addi
		disk[828] <= 32'b010010_11110_11011_1111111111111101; 	// sw
		disk[829] <= 32'b001111_11110_01010_1111111111111101; 	// lw
		disk[830] <= 32'b010110_00000000000000000000001001; 	// j
		disk[831] <= 32'b001110_01110_00001_0000000000000000; 	// mov
		disk[832] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[833] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[834] <= 32'b010000_00000_10100_0000000000001011; 	// li
		disk[835] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[836] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[837] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[838] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[839] <= 32'b010111_00000000000000000000000001; 	// jal
		disk[840] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[841] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[842] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[843] <= 32'b001110_01011_00110_0000000000000000; 	// mov
		disk[844] <= 32'b010000_00000_00111_0000000000000000; 	// li
		disk[845] <= 32'b010100_00000_00110_0000000000000000; 	// out
		disk[846] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[847] <= 32'b100101_11111_00000_0000000000000000; 	// syscall

		// PROGRAMA 2
		disk[850] <= 32'b010110_00000000000000000000011111;		// Jump to Main
		disk[851] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[852] <= 32'b010010_11110_00110_1111111111111100; 	// sw
		disk[853] <= 32'b010010_11110_00111_1111111111111101; 	// sw
		disk[854] <= 32'b010000_00000_10100_0000000000000000; 	// li
		disk[855] <= 32'b010010_11110_10100_1111111111111110; 	// sw
		disk[856] <= 32'b010000_00000_10101_0000000000000000; 	// li
		disk[857] <= 32'b010010_11110_10101_0000000000000000; 	// sw
		disk[858] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[859] <= 32'b001111_11110_01011_1111111111111101; 	// lw
		disk[860] <= 32'b000000_01010_01011_10110_00000_001110; 	// lt
		disk[861] <= 32'b010101_10110_00000_0000000000011011; 	// jf
		disk[862] <= 32'b001111_11110_01100_1111111111111100; 	// lw
		disk[863] <= 32'b000000_01100_01010_10111_00000_000000; 	// add
		disk[864] <= 32'b001111_10111_10111_0000000000000000; 	// lw
		disk[865] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[866] <= 32'b000000_01101_10111_11000_00000_001110; 	// lt
		disk[867] <= 32'b010101_11000_00000_0000000000010111; 	// jf
		disk[868] <= 32'b000000_01100_01010_11001_00000_000000; 	// add
		disk[869] <= 32'b001111_11001_11001_0000000000000000; 	// lw
		disk[870] <= 32'b010010_11110_11001_0000000000000000; 	// sw
		disk[871] <= 32'b001111_11110_01101_0000000000000000; 	// lw
		disk[872] <= 32'b010010_11110_01010_1111111111111111; 	// sw
		disk[873] <= 32'b000001_01010_11010_0000000000000001; 	// addi
		disk[874] <= 32'b010010_11110_11010_1111111111111110; 	// sw
		disk[875] <= 32'b001111_11110_01010_1111111111111110; 	// lw
		disk[876] <= 32'b010110_00000000000000000000001000; 	// j
		disk[877] <= 32'b001110_01101_00110_0000000000000000; 	// mov
		disk[878] <= 32'b010000_00000_00111_0000000000000001; 	// li
		disk[879] <= 32'b010100_00000_00110_0000000000000001; 	// out
		disk[880] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[881] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[882] <= 32'b010001_11110_01010_1111111111111011; 	// la
		disk[883] <= 32'b010000_00000_10100_0000000000001100; 	// li
		disk[884] <= 32'b010010_01010_10100_0000000000000000; 	// sw
		disk[885] <= 32'b010000_00000_10101_0000000000101001; 	// li
		disk[886] <= 32'b010010_01010_10101_0000000000000001; 	// sw
		disk[887] <= 32'b010000_00000_10110_0000000000010111; 	// li
		disk[888] <= 32'b010010_01010_10110_0000000000000010; 	// sw
		disk[889] <= 32'b010000_00000_10111_0000000001100010; 	// li
		disk[890] <= 32'b010010_01010_10111_0000000000000011; 	// sw
		disk[891] <= 32'b010000_00000_11000_0000000000100001; 	// li
		disk[892] <= 32'b010010_01010_11000_0000000000000100; 	// sw
		disk[893] <= 32'b010000_00000_11001_0000000000010101; 	// li
		disk[894] <= 32'b010010_01010_11001_0000000000000101; 	// sw
		disk[895] <= 32'b010001_11110_00110_1111111111111011; 	// la
		disk[896] <= 32'b010000_00000_00111_0000000000000110; 	// li
		disk[897] <= 32'b010010_11110_11111_1111111111111010; 	// sw
		disk[898] <= 32'b010111_00000000000000000000000001; 	// jal
		disk[899] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[900] <= 32'b001111_11110_11111_1111111111111010; 	// lw
		disk[901] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[902] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[903] <= 32'b100101_11111_00000_0000000000000000; 	// syscall
		
		// PROGRAMA 3
		disk[950] <= 32'b010110_00000000000000000000010011;		// Jump to Main
		disk[951] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[952] <= 32'b010010_11110_00110_1111111111111111; 	// sw
		disk[953] <= 32'b010000_00000_10100_0000000000000001; 	// li
		disk[954] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[955] <= 32'b001111_11110_01010_1111111111111111; 	// lw
		disk[956] <= 32'b010000_00000_10110_0000000000000000; 	// li
		disk[957] <= 32'b000000_01010_10110_10101_00000_010000; 	// gt
		disk[958] <= 32'b010101_10101_00000_0000000000010001; 	// jf
		disk[959] <= 32'b001111_11110_01011_0000000000000000; 	// lw
		disk[960] <= 32'b000000_01011_01010_10111_00000_000010; 	// mul
		disk[961] <= 32'b010010_11110_10111_0000000000000000; 	// sw
		disk[962] <= 32'b001111_11110_01011_0000000000000000; 	// lw
		disk[963] <= 32'b000010_01010_11000_0000000000000001; 	// subi
		disk[964] <= 32'b010010_11110_11000_1111111111111111; 	// sw
		disk[965] <= 32'b001111_11110_01010_1111111111111111; 	// lw
		disk[966] <= 32'b010110_00000000000000000000000101; 	// j
		disk[967] <= 32'b001110_01011_00001_0000000000000000; 	// mov
		disk[968] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[969] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[970] <= 32'b010000_00000_10100_0000000000000111; 	// li
		disk[971] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[972] <= 32'b001111_11110_01010_0000000000000000; 	// lw
		disk[973] <= 32'b001110_01010_00110_0000000000000000; 	// mov
		disk[974] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[975] <= 32'b010111_00000000000000000000000001; 	// jal
		disk[976] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[977] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[978] <= 32'b001110_00001_01011_0000000000000000; 	// mov
		disk[979] <= 32'b001110_01011_00110_0000000000000000; 	// mov
		disk[980] <= 32'b010000_00000_00111_0000000000000010; 	// li
		disk[981] <= 32'b010100_00000_00110_0000000000000010; 	// out
		disk[982] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[983] <= 32'b100101_11111_00000_0000000000000000; 	// syscall
		
	end
endmodule
