library verilog;
use verilog.vl_types.all;
entity iZero_vlg_vec_tst is
end iZero_vlg_vec_tst;
