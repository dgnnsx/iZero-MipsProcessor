module disco_rigido (clk, we, addr, datain, dataout);
	input clk;										// clock
	input we;										// write enable
	input [31:0] addr;							// disk address
	input [31:0] datain;							// data in (to disk)
	
	output reg [31:0] dataout;					// data out (from disk)
	
	localparam DISK_SIZE = 2048;				// Tamanho do disco
	reg [31:0] disk [DISK_SIZE-1:0];			// disk cells
	
	always @ (posedge clk) begin
		if (we) disk[addr] <= datain;			// write disk
	end
	
	always @ (negedge clk) begin
		dataout <= disk[addr];
	end

	initial begin
		// SISTEMA OPERACIONAL

disk[0] <= 32'b111100_00000000000000001001111110;		// Jump to Main
disk[1] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[2] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[3] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[4] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[5] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[6] <= 32'b010110_00001_10000_0000000000000000; 	// ldk
disk[7] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[8] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[9] <= 32'b001101_00101_10001_0000000000011010; 	// srli
disk[10] <= 32'b001111_11101_00110_0000000010100010; 	// lw
disk[11] <= 32'b000000_10001_00110_10010_00000_001101; 	// ne
disk[12] <= 32'b010101_10010_00000_0000000000010110; 	// jf
disk[13] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[14] <= 32'b000001_00111_10011_0000000000000001; 	// addi
disk[15] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[16] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[17] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[18] <= 32'b010110_00001_10100_0000000000000000; 	// ldk
disk[19] <= 32'b010010_11110_10100_1111111111111111; 	// sw
disk[20] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[21] <= 32'b111100_00000000000000000000001000; 	// j
disk[22] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[23] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[24] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[25] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[26] <= 32'b010010_11110_00001_1111111111111111; 	// sw
disk[27] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[28] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[29] <= 32'b000000_00101_10000_01111_00000_001100; 	// eq
disk[30] <= 32'b010101_01111_00000_0000000000100010; 	// jf
disk[31] <= 32'b010000_00000_10001_0000000000000001; 	// li
disk[32] <= 32'b001110_10001_11001_0000000000000000; 	// mov
disk[33] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[34] <= 32'b010000_00000_10010_0000000000000001; 	// li
disk[35] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[36] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[37] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[38] <= 32'b000000_00101_10100_10011_00000_010000; 	// gt
disk[39] <= 32'b010101_10011_00000_0000000000110000; 	// jf
disk[40] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[41] <= 32'b000011_00110_10101_0000000000000010; 	// muli
disk[42] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[43] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[44] <= 32'b000010_00101_10110_0000000000000001; 	// subi
disk[45] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[46] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[47] <= 32'b111100_00000000000000000000100100; 	// j
disk[48] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[49] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[50] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[51] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[52] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[53] <= 32'b010000_00000_00010_0000000000000000; 	// li
disk[54] <= 32'b010100_00000_00001_0000000000000000; 	// out
disk[55] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[56] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[57] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[58] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[59] <= 32'b010000_00000_00010_0000000000000010; 	// li
disk[60] <= 32'b010100_00000_00001_0000000000000010; 	// out
disk[61] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[62] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[63] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[64] <= 32'b010010_11101_01111_0000000001110011; 	// sw
disk[65] <= 32'b010000_00000_10000_0000000000000001; 	// li
disk[66] <= 32'b010010_11101_10000_0000000001110110; 	// sw
disk[67] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[68] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[69] <= 32'b010000_00000_01111_0000000000000001; 	// li
disk[70] <= 32'b010010_11101_01111_0000000000000000; 	// sw
disk[71] <= 32'b010000_00000_10000_0000000000000010; 	// li
disk[72] <= 32'b010010_11101_10000_0000000000000001; 	// sw
disk[73] <= 32'b010000_00000_10001_0000000000000011; 	// li
disk[74] <= 32'b010010_11101_10001_0000000000000010; 	// sw
disk[75] <= 32'b010000_00000_10010_0000000110010100; 	// li
disk[76] <= 32'b010010_11101_10010_0000000000000011; 	// sw
disk[77] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[78] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[79] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[80] <= 32'b010000_00000_10101_0000000000001010; 	// li
disk[81] <= 32'b000000_00101_10101_10100_00000_001110; 	// lt
disk[82] <= 32'b010101_10100_00000_0000000001100111; 	// jf
disk[83] <= 32'b010001_11101_00110_0000000000000100; 	// la
disk[84] <= 32'b000000_00110_00101_10110_00000_000000; 	// add
disk[85] <= 32'b010000_00000_10111_0000000000000000; 	// li
disk[86] <= 32'b010010_10110_10111_0000000000000000; 	// sw
disk[87] <= 32'b010001_11101_00111_0000000000001110; 	// la
disk[88] <= 32'b000000_00111_00101_11000_00000_000000; 	// add
disk[89] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[90] <= 32'b010010_11000_01111_0000000000000000; 	// sw
disk[91] <= 32'b010001_11101_01000_0000000000011000; 	// la
disk[92] <= 32'b000000_01000_00101_10000_00000_000000; 	// add
disk[93] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[94] <= 32'b010010_10000_10001_0000000000000000; 	// sw
disk[95] <= 32'b010001_11101_01001_0000000000100010; 	// la
disk[96] <= 32'b000000_01001_00101_10010_00000_000000; 	// add
disk[97] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[98] <= 32'b010010_10010_10011_0000000000000000; 	// sw
disk[99] <= 32'b000001_00101_10100_0000000000000001; 	// addi
disk[100] <= 32'b010010_11110_10100_0000000000000000; 	// sw
disk[101] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[102] <= 32'b111100_00000000000000000001001111; 	// j
disk[103] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[104] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[105] <= 32'b010000_00000_01111_0000000000100000; 	// li
disk[106] <= 32'b010010_11101_01111_0000000001101101; 	// sw
disk[107] <= 32'b010000_00000_10000_0000000001000000; 	// li
disk[108] <= 32'b010010_11101_10000_0000000001101110; 	// sw
disk[109] <= 32'b010000_00000_10001_0000000001100100; 	// li
disk[110] <= 32'b010010_11101_10001_0000000001101111; 	// sw
disk[111] <= 32'b010000_00000_10010_0000000000001010; 	// li
disk[112] <= 32'b010010_11101_10010_0000000001110000; 	// sw
disk[113] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[114] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[115] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[116] <= 32'b010010_11101_01111_0000000010100011; 	// sw
disk[117] <= 32'b010000_00000_10000_0000000000000001; 	// li
disk[118] <= 32'b010010_11101_10000_0000000010100100; 	// sw
disk[119] <= 32'b010000_00000_10001_0000000000000010; 	// li
disk[120] <= 32'b010010_11101_10001_0000000010100101; 	// sw
disk[121] <= 32'b010000_00000_10010_0000000000000011; 	// li
disk[122] <= 32'b010010_11101_10010_0000000010100110; 	// sw
disk[123] <= 32'b010000_00000_10011_0000000000000100; 	// li
disk[124] <= 32'b010010_11101_10011_0000000010100111; 	// sw
disk[125] <= 32'b010000_00000_10100_0000000000000101; 	// li
disk[126] <= 32'b010010_11101_10100_0000000010101000; 	// sw
disk[127] <= 32'b010000_00000_10101_0000000000001010; 	// li
disk[128] <= 32'b010010_11101_10101_0000000010101001; 	// sw
disk[129] <= 32'b001111_11101_00101_0000000010100011; 	// lw
disk[130] <= 32'b010010_11101_00101_0000000010101010; 	// sw
disk[131] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[132] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[133] <= 32'b010000_00000_01111_0000011111111111; 	// li
disk[134] <= 32'b010010_11101_01111_0000000001110010; 	// sw
disk[135] <= 32'b010000_00000_10000_0000000000011111; 	// li
disk[136] <= 32'b010010_11101_10000_0000000010100000; 	// sw
disk[137] <= 32'b010000_00000_10001_0000000000111101; 	// li
disk[138] <= 32'b010010_11101_10001_0000000010100001; 	// sw
disk[139] <= 32'b010000_00000_10010_0000000000111111; 	// li
disk[140] <= 32'b010010_11101_10010_0000000010100010; 	// sw
disk[141] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[142] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[143] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[144] <= 32'b010010_11110_01111_1111111111111110; 	// sw
disk[145] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[146] <= 32'b001111_11101_00110_0000000001101110; 	// lw
disk[147] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[148] <= 32'b010101_10000_00000_0000000010011101; 	// jf
disk[149] <= 32'b010001_11101_00111_0000000000101101; 	// la
disk[150] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[151] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[152] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[153] <= 32'b000001_00101_10011_0000000000000001; 	// addi
disk[154] <= 32'b010010_11110_10011_1111111111111110; 	// sw
disk[155] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[156] <= 32'b111100_00000000000000000010010001; 	// j
disk[157] <= 32'b010010_11110_11111_1111111111111101; 	// sw
disk[158] <= 32'b111110_00000000000000000000000001; 	// jal
disk[159] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[160] <= 32'b001111_11110_11111_1111111111111101; 	// lw
disk[161] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[162] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[163] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[164] <= 32'b000001_00110_10100_0000000000000001; 	// addi
disk[165] <= 32'b010010_11101_10100_0000000001110001; 	// sw
disk[166] <= 32'b001111_11101_00111_0000000001101101; 	// lw
disk[167] <= 32'b000000_00110_00111_10101_00000_000011; 	// div
disk[168] <= 32'b010010_11110_10101_1111111111111111; 	// sw
disk[169] <= 32'b000000_00110_00111_10110_00000_000100; 	// mod
disk[170] <= 32'b010000_00000_11000_0000000000000000; 	// li
disk[171] <= 32'b000000_10110_11000_10111_00000_010000; 	// gt
disk[172] <= 32'b010101_10111_00000_0000000010110001; 	// jf
disk[173] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[174] <= 32'b000001_01000_01111_0000000000000001; 	// addi
disk[175] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[176] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[177] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[178] <= 32'b010010_11110_10000_1111111111111110; 	// sw
disk[179] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[180] <= 32'b001111_11110_00110_1111111111111111; 	// lw
disk[181] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[182] <= 32'b010101_10001_00000_0000000010111111; 	// jf
disk[183] <= 32'b010001_11101_00111_0000000000101101; 	// la
disk[184] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
disk[185] <= 32'b010000_00000_10011_0000000000000001; 	// li
disk[186] <= 32'b010010_10010_10011_0000000000000000; 	// sw
disk[187] <= 32'b000001_00101_10100_0000000000000001; 	// addi
disk[188] <= 32'b010010_11110_10100_1111111111111110; 	// sw
disk[189] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[190] <= 32'b111100_00000000000000000010110011; 	// j
disk[191] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[192] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[193] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[194] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[195] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[196] <= 32'b001111_11101_00110_0000000001110000; 	// lw
disk[197] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[198] <= 32'b010101_10000_00000_0000000011011011; 	// jf
disk[199] <= 32'b010001_11101_00111_0000000001111000; 	// la
disk[200] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[201] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[202] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[203] <= 32'b010001_11101_01000_0000000010000010; 	// la
disk[204] <= 32'b000000_01000_00101_10011_00000_000000; 	// add
disk[205] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[206] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[207] <= 32'b010001_11101_01001_0000000010001100; 	// la
disk[208] <= 32'b000000_01001_00101_10101_00000_000000; 	// add
disk[209] <= 32'b010000_00000_10110_0000000000000000; 	// li
disk[210] <= 32'b010010_10101_10110_0000000000000000; 	// sw
disk[211] <= 32'b010001_11101_01010_0000000010010110; 	// la
disk[212] <= 32'b000000_01010_00101_10111_00000_000000; 	// add
disk[213] <= 32'b010000_00000_11000_0000000000000000; 	// li
disk[214] <= 32'b010010_10111_11000_0000000000000000; 	// sw
disk[215] <= 32'b000001_00101_01111_0000000000000001; 	// addi
disk[216] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[217] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[218] <= 32'b111100_00000000000000000011000011; 	// j
disk[219] <= 32'b001111_11101_00101_0000000001110001; 	// lw
disk[220] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[221] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[222] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[223] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[224] <= 32'b001111_11101_00110_0000000001110010; 	// lw
disk[225] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[226] <= 32'b010101_10001_00000_0000000011111011; 	// jf
disk[227] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[228] <= 32'b010110_00001_10010_0000000000000000; 	// ldk
disk[229] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[230] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[231] <= 32'b001101_00111_10011_0000000000011010; 	// srli
disk[232] <= 32'b001111_11101_01000_0000000010100001; 	// lw
disk[233] <= 32'b000000_10011_01000_10100_00000_001100; 	// eq
disk[234] <= 32'b010101_10100_00000_0000000011110110; 	// jf
disk[235] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[236] <= 32'b000001_01001_10101_0000000000000001; 	// addi
disk[237] <= 32'b010001_11101_01010_0000000001111000; 	// la
disk[238] <= 32'b000000_01010_01001_10110_00000_000000; 	// add
disk[239] <= 32'b010010_10110_10101_0000000000000000; 	// sw
disk[240] <= 32'b010001_11101_01011_0000000010000010; 	// la
disk[241] <= 32'b000000_01011_01001_10111_00000_000000; 	// add
disk[242] <= 32'b010010_10111_00101_0000000000000000; 	// sw
disk[243] <= 32'b000001_01001_11000_0000000000000001; 	// addi
disk[244] <= 32'b010010_11110_11000_1111111111111111; 	// sw
disk[245] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[246] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[247] <= 32'b000001_00101_01111_0000000000000001; 	// addi
disk[248] <= 32'b010010_11110_01111_1111111111111110; 	// sw
disk[249] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[250] <= 32'b111100_00000000000000000011011111; 	// j
disk[251] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[252] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[253] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[254] <= 32'b111110_00000000000000000001000100; 	// jal
disk[255] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[256] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[257] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[258] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[259] <= 32'b111110_00000000000000000001101000; 	// jal
disk[260] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[261] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[262] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[263] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[264] <= 32'b111110_00000000000000000001110010; 	// jal
disk[265] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[266] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[267] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[268] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[269] <= 32'b111110_00000000000000000010000100; 	// jal
disk[270] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[271] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[272] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[273] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[274] <= 32'b111110_00000000000000000010001110; 	// jal
disk[275] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[276] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[277] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[278] <= 32'b010010_11110_11111_0000000000000000; 	// sw
disk[279] <= 32'b111110_00000000000000000011000000; 	// jal
disk[280] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[281] <= 32'b001111_11110_11111_0000000000000000; 	// lw
disk[282] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[283] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[284] <= 32'b000001_11110_11110_0000000000000110; 	// addi
disk[285] <= 32'b010010_11110_00001_1111111111111101; 	// sw
disk[286] <= 32'b001111_11110_00101_1111111111111101; 	// lw
disk[287] <= 32'b001111_11101_00110_0000000001101101; 	// lw
disk[288] <= 32'b000000_00101_00110_01111_00000_000011; 	// div
disk[289] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[290] <= 32'b000000_00101_00110_10000_00000_000100; 	// mod
disk[291] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[292] <= 32'b000000_10000_10010_10001_00000_010000; 	// gt
disk[293] <= 32'b010101_10001_00000_0000000100101010; 	// jf
disk[294] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[295] <= 32'b000001_00111_10011_0000000000000001; 	// addi
disk[296] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[297] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[298] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[299] <= 32'b010010_11110_10100_1111111111111110; 	// sw
disk[300] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[301] <= 32'b001111_11101_00110_0000000001101110; 	// lw
disk[302] <= 32'b000000_00101_00110_10101_00000_001110; 	// lt
disk[303] <= 32'b010101_10101_00000_0000000101001111; 	// jf
disk[304] <= 32'b010001_11101_00111_0000000000101101; 	// la
disk[305] <= 32'b000000_00111_00101_10110_00000_000000; 	// add
disk[306] <= 32'b001111_10110_10110_0000000000000000; 	// lw
disk[307] <= 32'b010000_00000_11000_0000000000000000; 	// li
disk[308] <= 32'b000000_10110_11000_10111_00000_001100; 	// eq
disk[309] <= 32'b010101_10111_00000_0000000101001010; 	// jf
disk[310] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[311] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[312] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[313] <= 32'b000000_00101_10000_01111_00000_001101; 	// ne
disk[314] <= 32'b010101_01111_00000_0000000101000111; 	// jf
disk[315] <= 32'b010001_11101_00110_0000000000101101; 	// la
disk[316] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[317] <= 32'b000000_00110_00111_10001_00000_000000; 	// add
disk[318] <= 32'b010000_00000_10010_0000000000000001; 	// li
disk[319] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[320] <= 32'b000010_00101_10011_0000000000000001; 	// subi
disk[321] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[322] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[323] <= 32'b000001_00111_10100_0000000000000001; 	// addi
disk[324] <= 32'b010010_11110_10100_1111111111111110; 	// sw
disk[325] <= 32'b001111_11110_00111_1111111111111110; 	// lw
disk[326] <= 32'b111100_00000000000000000100110111; 	// j
disk[327] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[328] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[329] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[330] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[331] <= 32'b000001_00101_10101_0000000000000001; 	// addi
disk[332] <= 32'b010010_11110_10101_1111111111111110; 	// sw
disk[333] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[334] <= 32'b111100_00000000000000000100101100; 	// j
disk[335] <= 32'b001111_11101_00101_0000000001101111; 	// lw
disk[336] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[337] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[338] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[339] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[340] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[341] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[342] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[343] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[344] <= 32'b001111_11101_00110_0000000001110000; 	// lw
disk[345] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[346] <= 32'b010101_10001_00000_0000000101110000; 	// jf
disk[347] <= 32'b010001_11101_00111_0000000010001100; 	// la
disk[348] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
disk[349] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[350] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[351] <= 32'b000000_10010_10100_10011_00000_001101; 	// ne
disk[352] <= 32'b010101_10011_00000_0000000101101011; 	// jf
disk[353] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[354] <= 32'b010010_11110_11111_1111111111111110; 	// sw
disk[355] <= 32'b111110_00000000000000000000011001; 	// jal
disk[356] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[357] <= 32'b001111_11110_11111_1111111111111110; 	// lw
disk[358] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[359] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[360] <= 32'b000000_00110_00101_10101_00000_000000; 	// add
disk[361] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[362] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[363] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[364] <= 32'b000001_00101_10110_0000000000000001; 	// addi
disk[365] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[366] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[367] <= 32'b111100_00000000000000000101010111; 	// j
disk[368] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[369] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[370] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[371] <= 32'b000001_11110_11110_0000000000000100; 	// addi
disk[372] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[373] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[374] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[375] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[376] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[377] <= 32'b001111_11101_00110_0000000001110000; 	// lw
disk[378] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
disk[379] <= 32'b010101_10001_00000_0000000110010001; 	// jf
disk[380] <= 32'b010001_11101_00111_0000000001111000; 	// la
disk[381] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
disk[382] <= 32'b001111_10010_10010_0000000000000000; 	// lw
disk[383] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[384] <= 32'b000000_10010_10100_10011_00000_001101; 	// ne
disk[385] <= 32'b010101_10011_00000_0000000110001100; 	// jf
disk[386] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[387] <= 32'b010010_11110_11111_1111111111111110; 	// sw
disk[388] <= 32'b111110_00000000000000000000011001; 	// jal
disk[389] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[390] <= 32'b001111_11110_11111_1111111111111110; 	// lw
disk[391] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[392] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[393] <= 32'b000000_00110_00101_10101_00000_000000; 	// add
disk[394] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[395] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[396] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[397] <= 32'b000001_00101_10110_0000000000000001; 	// addi
disk[398] <= 32'b010010_11110_10110_1111111111111111; 	// sw
disk[399] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[400] <= 32'b111100_00000000000000000101111000; 	// j
disk[401] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[402] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[403] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[404] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[405] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[406] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[407] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[408] <= 32'b001111_11101_00110_0000000001110000; 	// lw
disk[409] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[410] <= 32'b010101_10000_00000_0000000110101000; 	// jf
disk[411] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[412] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[413] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[414] <= 32'b001111_11101_01000_0000000000000010; 	// lw
disk[415] <= 32'b000000_10001_01000_10010_00000_001100; 	// eq
disk[416] <= 32'b010101_10010_00000_0000000110100011; 	// jf
disk[417] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[418] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[419] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[420] <= 32'b000001_00101_10011_0000000000000001; 	// addi
disk[421] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[422] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[423] <= 32'b111100_00000000000000000110010111; 	// j
disk[424] <= 32'b001111_11101_00101_0000000000000011; 	// lw
disk[425] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[426] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[427] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[428] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[429] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[430] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[431] <= 32'b001111_11101_00110_0000000001110000; 	// lw
disk[432] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[433] <= 32'b010101_10000_00000_0000000110111111; 	// jf
disk[434] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[435] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[436] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[437] <= 32'b001111_11101_01000_0000000000000001; 	// lw
disk[438] <= 32'b000000_10001_01000_10010_00000_001100; 	// eq
disk[439] <= 32'b010101_10010_00000_0000000110111010; 	// jf
disk[440] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[441] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[442] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[443] <= 32'b000001_00101_10011_0000000000000001; 	// addi
disk[444] <= 32'b010010_11110_10011_0000000000000000; 	// sw
disk[445] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[446] <= 32'b111100_00000000000000000110101110; 	// j
disk[447] <= 32'b001111_11101_00101_0000000000000011; 	// lw
disk[448] <= 32'b001110_00101_11001_0000000000000000; 	// mov
disk[449] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[450] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[451] <= 32'b010000_00000_01111_0000000000000000; 	// li
disk[452] <= 32'b010010_11110_01111_0000000000000000; 	// sw
disk[453] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[454] <= 32'b001111_11101_00110_0000000001110000; 	// lw
disk[455] <= 32'b000000_00101_00110_10000_00000_001110; 	// lt
disk[456] <= 32'b010101_10000_00000_0000000111011000; 	// jf
disk[457] <= 32'b010001_11101_00111_0000000010001100; 	// la
disk[458] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[459] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[460] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[461] <= 32'b000000_10001_10011_10010_00000_001101; 	// ne
disk[462] <= 32'b010101_10010_00000_0000000111010011; 	// jf
disk[463] <= 32'b010001_11101_01000_0000000000000100; 	// la
disk[464] <= 32'b000000_01000_00101_10100_00000_000000; 	// add
disk[465] <= 32'b001111_11101_01001_0000000000000001; 	// lw
disk[466] <= 32'b010010_10100_01001_0000000000000000; 	// sw
disk[467] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[468] <= 32'b000001_00101_10101_0000000000000001; 	// addi
disk[469] <= 32'b010010_11110_10101_0000000000000000; 	// sw
disk[470] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[471] <= 32'b111100_00000000000000000111000101; 	// j
disk[472] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[473] <= 32'b000001_11110_11110_0000000000000101; 	// addi
disk[474] <= 32'b010010_11110_00001_1111111111111110; 	// sw
disk[475] <= 32'b001111_11110_00101_1111111111111110; 	// lw
disk[476] <= 32'b010010_11110_00101_0000000000000000; 	// sw
disk[477] <= 32'b001111_11110_00110_0000000000000000; 	// lw
disk[478] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[479] <= 32'b010110_00001_01111_0000000000000000; 	// ldk
disk[480] <= 32'b010010_11110_01111_1111111111111111; 	// sw
disk[481] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[482] <= 32'b001101_00101_10000_0000000000011010; 	// srli
disk[483] <= 32'b001111_11101_00110_0000000010100000; 	// lw
disk[484] <= 32'b000000_10000_00110_10001_00000_001101; 	// ne
disk[485] <= 32'b010101_10001_00000_0000000111101111; 	// jf
disk[486] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[487] <= 32'b000001_00111_10010_0000000000000001; 	// addi
disk[488] <= 32'b010010_11110_10010_0000000000000000; 	// sw
disk[489] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[490] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[491] <= 32'b010110_00001_10011_0000000000000000; 	// ldk
disk[492] <= 32'b010010_11110_10011_1111111111111111; 	// sw
disk[493] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[494] <= 32'b111100_00000000000000000111100001; 	// j
disk[495] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[496] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[497] <= 32'b000000_00101_00110_10100_00000_000001; 	// sub
disk[498] <= 32'b001110_10100_11001_0000000000000000; 	// mov
disk[499] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[500] <= 32'b000001_11110_11110_0000000000001010; 	// addi
disk[501] <= 32'b010010_11110_00001_1111111111111001; 	// sw
disk[502] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[503] <= 32'b000010_00101_01111_0000000000000001; 	// subi
disk[504] <= 32'b010010_11110_01111_1111111111111001; 	// sw
disk[505] <= 32'b001111_11110_00101_1111111111111001; 	// lw
disk[506] <= 32'b010001_11101_00110_0000000010000010; 	// la
disk[507] <= 32'b000000_00110_00101_10000_00000_000000; 	// add
disk[508] <= 32'b001111_10000_10000_0000000000000000; 	// lw
disk[509] <= 32'b010010_11110_10000_1111111111111111; 	// sw
disk[510] <= 32'b010001_11101_00111_0000000001111000; 	// la
disk[511] <= 32'b000000_00111_00101_10001_00000_000000; 	// add
disk[512] <= 32'b001111_10001_10001_0000000000000000; 	// lw
disk[513] <= 32'b010010_11110_10001_0000000000000000; 	// sw
disk[514] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[515] <= 32'b010010_11110_01000_1111111111111010; 	// sw
disk[516] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[517] <= 32'b010010_11110_11111_1111111111111000; 	// sw
disk[518] <= 32'b111110_00000000000000000111011001; 	// jal
disk[519] <= 32'b000010_11110_11110_0000000000000101; 	// subi
disk[520] <= 32'b001111_11110_11111_1111111111111000; 	// lw
disk[521] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[522] <= 32'b010010_11110_00101_1111111111111110; 	// sw
disk[523] <= 32'b001111_11110_00110_1111111111111110; 	// lw
disk[524] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[525] <= 32'b010010_11110_11111_1111111111111000; 	// sw
disk[526] <= 32'b111110_00000000000000000100011100; 	// jal
disk[527] <= 32'b000010_11110_11110_0000000000000110; 	// subi
disk[528] <= 32'b001111_11110_11111_1111111111111000; 	// lw
disk[529] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[530] <= 32'b010010_11110_00101_1111111111111101; 	// sw
disk[531] <= 32'b001111_11101_00110_0000000001101101; 	// lw
disk[532] <= 32'b001111_11110_00111_1111111111111101; 	// lw
disk[533] <= 32'b000000_00110_00111_10010_00000_000010; 	// mul
disk[534] <= 32'b010010_11110_10010_1111111111111011; 	// sw
disk[535] <= 32'b001111_11110_01000_1111111111111010; 	// lw
disk[536] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[537] <= 32'b010110_00001_10011_0000000000000000; 	// ldk
disk[538] <= 32'b010010_11110_10011_1111111111111100; 	// sw
disk[539] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[540] <= 32'b001101_00101_10100_0000000000011010; 	// srli
disk[541] <= 32'b001111_11101_00110_0000000010100000; 	// lw
disk[542] <= 32'b000000_10100_00110_10101_00000_001101; 	// ne
disk[543] <= 32'b010101_10101_00000_0000001000110000; 	// jf
disk[544] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[545] <= 32'b001111_11110_00111_1111111111111011; 	// lw
disk[546] <= 32'b001110_00111_00010_0000000000000000; 	// mov
disk[547] <= 32'b011001_00010_00001_0000000000000000; 	// sim
disk[548] <= 32'b001111_11110_01000_1111111111111010; 	// lw
disk[549] <= 32'b000001_01000_10110_0000000000000001; 	// addi
disk[550] <= 32'b010010_11110_10110_1111111111111010; 	// sw
disk[551] <= 32'b001111_11110_01000_1111111111111010; 	// lw
disk[552] <= 32'b001110_01000_00001_0000000000000000; 	// mov
disk[553] <= 32'b010110_00001_10111_0000000000000000; 	// ldk
disk[554] <= 32'b010010_11110_10111_1111111111111100; 	// sw
disk[555] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[556] <= 32'b000001_00111_11000_0000000000000001; 	// addi
disk[557] <= 32'b010010_11110_11000_1111111111111011; 	// sw
disk[558] <= 32'b001111_11110_00111_1111111111111011; 	// lw
disk[559] <= 32'b111100_00000000000000001000011011; 	// j
disk[560] <= 32'b001111_11110_00101_1111111111111100; 	// lw
disk[561] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[562] <= 32'b001111_11110_00110_1111111111111011; 	// lw
disk[563] <= 32'b001110_00110_00010_0000000000000000; 	// mov
disk[564] <= 32'b011001_00010_00001_0000000000000000; 	// sim
disk[565] <= 32'b001111_11110_00111_0000000000000000; 	// lw
disk[566] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[567] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
disk[568] <= 32'b001111_11101_01000_0000000001101101; 	// lw
disk[569] <= 32'b001111_11110_01001_1111111111111101; 	// lw
disk[570] <= 32'b000000_01000_01001_01111_00000_000010; 	// mul
disk[571] <= 32'b001110_01111_00001_0000000000000000; 	// mov
disk[572] <= 32'b011010_00000_00001_0000000000000000; 	// mmuLowerIM
disk[573] <= 32'b010001_11101_01010_0000000010001100; 	// la
disk[574] <= 32'b001111_11110_01011_1111111111111001; 	// lw
disk[575] <= 32'b000000_01010_01011_10000_00000_000000; 	// add
disk[576] <= 32'b010010_10000_00111_0000000000000000; 	// sw
disk[577] <= 32'b010001_11101_01100_0000000010010110; 	// la
disk[578] <= 32'b000000_01100_01011_10001_00000_000000; 	// add
disk[579] <= 32'b001111_11110_01101_1111111111111111; 	// lw
disk[580] <= 32'b010010_10001_01101_0000000000000000; 	// sw
disk[581] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[582] <= 32'b000001_11110_11110_0000000000000011; 	// addi
disk[583] <= 32'b010010_11110_00001_0000000000000000; 	// sw
disk[584] <= 32'b001111_11110_00101_0000000000000000; 	// lw
disk[585] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[586] <= 32'b100100_00000_00001_0000000000000000; 	// lcdCurr
disk[587] <= 32'b001111_11101_00110_0000000010101001; 	// lw
disk[588] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[589] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[590] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[591] <= 32'b001111_11101_01000_0000000000101100; 	// lw
disk[592] <= 32'b000000_00111_01000_01111_00000_000000; 	// add
disk[593] <= 32'b001111_11101_01001_0000000000000000; 	// lw
disk[594] <= 32'b010010_01111_01001_0000000000000000; 	// sw
disk[595] <= 32'b010001_11101_01010_0000000000001110; 	// la
disk[596] <= 32'b000000_01010_01000_10000_00000_000000; 	// add
disk[597] <= 32'b010000_00000_10001_0000000000000000; 	// li
disk[598] <= 32'b010010_10000_10001_0000000000000000; 	// sw
disk[599] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[600] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
disk[601] <= 32'b010010_11110_11111_1111111111111111; 	// sw
disk[602] <= 32'b100000_00000000000000000000000000; 	// exec
disk[603] <= 32'b001111_11110_11111_1111111111111111; 	// lw
disk[604] <= 32'b000000_00111_01000_10010_00000_000000; 	// add
disk[605] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[606] <= 32'b010010_10010_10011_0000000000000000; 	// sw
disk[607] <= 32'b000000_01010_01000_10100_00000_000000; 	// add
disk[608] <= 32'b010000_00000_10101_0000000000000000; 	// li
disk[609] <= 32'b010010_10100_10101_0000000000000000; 	// sw
disk[610] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[611] <= 32'b000001_11110_11110_0000000000000010; 	// addi
disk[612] <= 32'b010010_11110_00001_0000000000000001; 	// sw
disk[613] <= 32'b001111_11110_00101_0000000000000001; 	// lw
disk[614] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[615] <= 32'b100100_00000_00001_0000000000000000; 	// lcdCurr
disk[616] <= 32'b001111_11101_00110_0000000010101001; 	// lw
disk[617] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[618] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[619] <= 32'b010001_11101_00111_0000000000000100; 	// la
disk[620] <= 32'b001111_11101_01000_0000000000101100; 	// lw
disk[621] <= 32'b000000_00111_01000_01111_00000_000000; 	// add
disk[622] <= 32'b001111_11101_01001_0000000000000000; 	// lw
disk[623] <= 32'b010010_01111_01001_0000000000000000; 	// sw
disk[624] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[625] <= 32'b010001_11101_01010_0000000000001110; 	// la
disk[626] <= 32'b000000_01010_01000_10000_00000_000000; 	// add
disk[627] <= 32'b001111_10000_10000_0000000000000000; 	// lw
disk[628] <= 32'b001110_10000_00010_0000000000000000; 	// mov
disk[629] <= 32'b011110_00001_00000_0000000000000000; 	// mmuSelect
disk[630] <= 32'b100001_00010_00000_0000000000000000; 	// execAgain
disk[631] <= 32'b000000_00111_01000_10001_00000_000000; 	// add
disk[632] <= 32'b010000_00000_10010_0000000000000000; 	// li
disk[633] <= 32'b010010_10001_10010_0000000000000000; 	// sw
disk[634] <= 32'b000000_01010_01000_10011_00000_000000; 	// add
disk[635] <= 32'b010000_00000_10100_0000000000000000; 	// li
disk[636] <= 32'b010010_10011_10100_0000000000000000; 	// sw
disk[637] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
disk[638] <= 32'b010000_00000_00000_0000000000000000; 	// li
disk[639] <= 32'b010000_00000_11110_0000000000000000; 	// li
disk[640] <= 32'b010000_00000_11101_0000000000000000; 	// li
disk[641] <= 32'b000001_11110_11110_0000000010101110; 	// addi
disk[642] <= 32'b111110_00000000000000000011111100; 	// jal
disk[643] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[644] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[645] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[646] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[647] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[648] <= 32'b010000_00000_00001_0000000000000000; 	// li
disk[649] <= 32'b001110_00001_11010_0000000000000000; 	// mov
disk[650] <= 32'b010000_00000_01111_0000000000000001; 	// li
disk[651] <= 32'b010101_01111_00000_0000001101010001; 	// jf
disk[652] <= 32'b001110_11010_10000_0000000000000000; 	// mov
disk[653] <= 32'b010010_11110_10000_0000000000000000; 	// sw
disk[654] <= 32'b010011_00000_10001_0000000000000000; 	// in
disk[655] <= 32'b010010_11110_10001_1111111111111111; 	// sw
disk[656] <= 32'b111110_00000000000000000101110011; 	// jal
disk[657] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[658] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[659] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[660] <= 32'b010000_00000_00010_0000000000000000; 	// li
disk[661] <= 32'b010100_00000_00001_0000000000000000; 	// out
disk[662] <= 32'b001111_11101_00110_0000000010101010; 	// lw
disk[663] <= 32'b001111_11101_00111_0000000010100011; 	// lw
disk[664] <= 32'b000000_00110_00111_10010_00000_001100; 	// eq
disk[665] <= 32'b010101_10010_00000_0000001010110011; 	// jf
disk[666] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[667] <= 32'b010000_00000_10100_0000000000000100; 	// li
disk[668] <= 32'b000000_01000_10100_10011_00000_010000; 	// gt
disk[669] <= 32'b010101_10011_00000_0000001010100001; 	// jf
disk[670] <= 32'b010010_11110_00111_1111111111111111; 	// sw
disk[671] <= 32'b001111_11110_01000_1111111111111111; 	// lw
disk[672] <= 32'b111100_00000000000000001010110010; 	// j
disk[673] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[674] <= 32'b010000_00000_10110_0000000000000100; 	// li
disk[675] <= 32'b000000_00101_10110_10101_00000_001100; 	// eq
disk[676] <= 32'b010101_10101_00000_0000001010101011; 	// jf
disk[677] <= 32'b111110_00000000000000000000110011; 	// jal
disk[678] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[679] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[680] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[681] <= 32'b010010_11110_00110_1111111111111111; 	// sw
disk[682] <= 32'b111100_00000000000000001010110010; 	// j
disk[683] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[684] <= 32'b010000_00000_11000_0000000000000001; 	// li
disk[685] <= 32'b000000_00101_11000_10111_00000_001110; 	// lt
disk[686] <= 32'b010101_10111_00000_0000001010110010; 	// jf
disk[687] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[688] <= 32'b010010_11110_00110_1111111111111111; 	// sw
disk[689] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[690] <= 32'b111100_00000000000000001101001011; 	// j
disk[691] <= 32'b001111_11101_00101_0000000010101010; 	// lw
disk[692] <= 32'b001111_11101_00110_0000000010100100; 	// lw
disk[693] <= 32'b000000_00101_00110_01111_00000_001100; 	// eq
disk[694] <= 32'b010101_01111_00000_0000001011000111; 	// jf
disk[695] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[696] <= 32'b010000_00000_10001_0000000000000011; 	// li
disk[697] <= 32'b000000_00111_10001_10000_00000_010000; 	// gt
disk[698] <= 32'b010101_10000_00000_0000001010111111; 	// jf
disk[699] <= 32'b001111_11101_01000_0000000010100011; 	// lw
disk[700] <= 32'b010010_11110_01000_1111111111111111; 	// sw
disk[701] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[702] <= 32'b111100_00000000000000001011000110; 	// j
disk[703] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[704] <= 32'b010000_00000_10011_0000000000000001; 	// li
disk[705] <= 32'b000000_00101_10011_10010_00000_001110; 	// lt
disk[706] <= 32'b010101_10010_00000_0000001011000110; 	// jf
disk[707] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[708] <= 32'b010010_11110_00110_1111111111111111; 	// sw
disk[709] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[710] <= 32'b111100_00000000000000001101001011; 	// j
disk[711] <= 32'b001111_11101_00101_0000000010101010; 	// lw
disk[712] <= 32'b001111_11101_00110_0000000010100101; 	// lw
disk[713] <= 32'b000000_00101_00110_10100_00000_001100; 	// eq
disk[714] <= 32'b010101_10100_00000_0000001011101000; 	// jf
disk[715] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[716] <= 32'b010000_00000_10110_0000000000000001; 	// li
disk[717] <= 32'b000000_00111_10110_10101_00000_001100; 	// eq
disk[718] <= 32'b010101_10101_00000_0000001011011000; 	// jf
disk[719] <= 32'b001111_11101_01000_0000000010100111; 	// lw
disk[720] <= 32'b010010_11110_01000_1111111111111111; 	// sw
disk[721] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[722] <= 32'b111110_00000000000000000101110011; 	// jal
disk[723] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[724] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[725] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[726] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[727] <= 32'b111100_00000000000000001011100111; 	// j
disk[728] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[729] <= 32'b010000_00000_11000_0000000000000011; 	// li
disk[730] <= 32'b000000_00101_11000_10111_00000_010000; 	// gt
disk[731] <= 32'b010101_10111_00000_0000001011100000; 	// jf
disk[732] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[733] <= 32'b010010_11110_00110_1111111111111111; 	// sw
disk[734] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[735] <= 32'b111100_00000000000000001011100111; 	// j
disk[736] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[737] <= 32'b010000_00000_10000_0000000000000001; 	// li
disk[738] <= 32'b000000_00101_10000_01111_00000_001110; 	// lt
disk[739] <= 32'b010101_01111_00000_0000001011100111; 	// jf
disk[740] <= 32'b001111_11101_00110_0000000010100011; 	// lw
disk[741] <= 32'b010010_11110_00110_1111111111111111; 	// sw
disk[742] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[743] <= 32'b111100_00000000000000001101001011; 	// j
disk[744] <= 32'b001111_11101_00101_0000000010101010; 	// lw
disk[745] <= 32'b001111_11101_00110_0000000010100110; 	// lw
disk[746] <= 32'b000000_00101_00110_10001_00000_001100; 	// eq
disk[747] <= 32'b010101_10001_00000_0000001100010110; 	// jf
disk[748] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[749] <= 32'b010000_00000_10011_0000000000000001; 	// li
disk[750] <= 32'b000000_00111_10011_10010_00000_001100; 	// eq
disk[751] <= 32'b010101_10010_00000_0000001100000111; 	// jf
disk[752] <= 32'b111110_00000000000000000111000010; 	// jal
disk[753] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[754] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[755] <= 32'b111110_00000000000000000110101011; 	// jal
disk[756] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[757] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[758] <= 32'b001111_11101_00110_0000000000000011; 	// lw
disk[759] <= 32'b000000_00101_00110_10100_00000_001101; 	// ne
disk[760] <= 32'b010101_10100_00000_0000001100000100; 	// jf
disk[761] <= 32'b111110_00000000000000000110101011; 	// jal
disk[762] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[763] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[764] <= 32'b010010_11101_00101_0000000000101100; 	// sw
disk[765] <= 32'b001111_11101_00110_0000000000101100; 	// lw
disk[766] <= 32'b000001_00110_10101_0000000000000001; 	// addi
disk[767] <= 32'b001110_10101_00001_0000000000000000; 	// mov
disk[768] <= 32'b111110_00000000000000001001000110; 	// jal
disk[769] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[770] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[771] <= 32'b111100_00000000000000001011110011; 	// j
disk[772] <= 32'b001111_11101_00101_0000000010100011; 	// lw
disk[773] <= 32'b010010_11110_00101_1111111111111111; 	// sw
disk[774] <= 32'b111100_00000000000000001100010101; 	// j
disk[775] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[776] <= 32'b010000_00000_10111_0000000000000010; 	// li
disk[777] <= 32'b000000_00101_10111_10110_00000_001100; 	// eq
disk[778] <= 32'b010101_10110_00000_0000001100010011; 	// jf
disk[779] <= 32'b111110_00000000000000000101010010; 	// jal
disk[780] <= 32'b000010_11110_11110_0000000000000100; 	// subi
disk[781] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[782] <= 32'b001110_00101_00001_0000000000000000; 	// mov
disk[783] <= 32'b100011_00000_00001_0000000000000000; 	// lcdPgms
disk[784] <= 32'b001111_11101_00110_0000000010101000; 	// lw
disk[785] <= 32'b010010_11110_00110_1111111111111111; 	// sw
disk[786] <= 32'b111100_00000000000000001100010101; 	// j
disk[787] <= 32'b001111_11101_00101_0000000010100011; 	// lw
disk[788] <= 32'b010010_11110_00101_1111111111111111; 	// sw
disk[789] <= 32'b111100_00000000000000001101001011; 	// j
disk[790] <= 32'b001111_11101_00101_0000000010101010; 	// lw
disk[791] <= 32'b001111_11101_00110_0000000010100111; 	// lw
disk[792] <= 32'b000000_00101_00110_11000_00000_001100; 	// eq
disk[793] <= 32'b010101_11000_00000_0000001100100101; 	// jf
disk[794] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[795] <= 32'b010000_00000_10000_0000000000000000; 	// li
disk[796] <= 32'b000000_00111_10000_01111_00000_010000; 	// gt
disk[797] <= 32'b010101_01111_00000_0000001100100010; 	// jf
disk[798] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[799] <= 32'b111110_00000000000000000111110100; 	// jal
disk[800] <= 32'b000010_11110_11110_0000000000001010; 	// subi
disk[801] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[802] <= 32'b001111_11101_00101_0000000010100011; 	// lw
disk[803] <= 32'b010010_11110_00101_1111111111111111; 	// sw
disk[804] <= 32'b111100_00000000000000001101001011; 	// j
disk[805] <= 32'b001111_11101_00101_0000000010101010; 	// lw
disk[806] <= 32'b001111_11101_00110_0000000010101000; 	// lw
disk[807] <= 32'b000000_00101_00110_10001_00000_001100; 	// eq
disk[808] <= 32'b010101_10001_00000_0000001101001011; 	// jf
disk[809] <= 32'b001111_11110_00111_1111111111111111; 	// lw
disk[810] <= 32'b010000_00000_10011_0000000000000000; 	// li
disk[811] <= 32'b000000_00111_10011_10010_00000_010000; 	// gt
disk[812] <= 32'b010101_10010_00000_0000001101001001; 	// jf
disk[813] <= 32'b000010_00111_10100_0000000000000001; 	// subi
disk[814] <= 32'b010010_11101_10100_0000000000101100; 	// sw
disk[815] <= 32'b001110_00111_00001_0000000000000000; 	// mov
disk[816] <= 32'b111110_00000000000000001001000110; 	// jal
disk[817] <= 32'b000010_11110_11110_0000000000000011; 	// subi
disk[818] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[819] <= 32'b010001_11101_00101_0000000000000100; 	// la
disk[820] <= 32'b001111_11101_00110_0000000000101100; 	// lw
disk[821] <= 32'b000000_00101_00110_10101_00000_000000; 	// add
disk[822] <= 32'b001111_10101_10101_0000000000000000; 	// lw
disk[823] <= 32'b001111_11101_00111_0000000000000010; 	// lw
disk[824] <= 32'b000000_10101_00111_10110_00000_001100; 	// eq
disk[825] <= 32'b010101_10110_00000_0000001101001001; 	// jf
disk[826] <= 32'b010001_11101_01000_0000000000001110; 	// la
disk[827] <= 32'b000000_01000_00110_10111_00000_000000; 	// add
disk[828] <= 32'b001111_10111_10111_0000000000000000; 	// lw
disk[829] <= 32'b001110_10111_00001_0000000000000000; 	// mov
disk[830] <= 32'b010000_00000_00010_0000000000000010; 	// li
disk[831] <= 32'b010100_00000_00001_0000000000000010; 	// out
disk[832] <= 32'b010000_00000_00001_0000000000100000; 	// li
disk[833] <= 32'b010000_00000_00010_0000000000000001; 	// li
disk[834] <= 32'b010100_00000_00001_0000000000000001; 	// out
disk[835] <= 32'b001111_11110_01001_1111111111111111; 	// lw
disk[836] <= 32'b001110_01001_00001_0000000000000000; 	// mov
disk[837] <= 32'b111110_00000000000000001001100011; 	// jal
disk[838] <= 32'b000010_11110_11110_0000000000000010; 	// subi
disk[839] <= 32'b001110_11001_00101_0000000000000000; 	// mov
disk[840] <= 32'b111100_00000000000000001100110011; 	// j
disk[841] <= 32'b001111_11101_00101_0000000010100011; 	// lw
disk[842] <= 32'b010010_11110_00101_1111111111111111; 	// sw
disk[843] <= 32'b001111_11110_00101_1111111111111111; 	// lw
disk[844] <= 32'b010010_11101_00101_0000000010101010; 	// sw
disk[845] <= 32'b001111_11101_00110_0000000010101010; 	// lw
disk[846] <= 32'b001110_00110_00001_0000000000000000; 	// mov
disk[847] <= 32'b100010_00000_00001_0000000000000000; 	// lcd
disk[848] <= 32'b111100_00000000000000001010001010; 	// j
disk[849] <= 32'b111111_00000000000000000000000000; 	// halt



		// PROGRAMA 1
		disk[1700] <= 32'b111101_00000000000000000000100011;		// Jump to Main
		disk[1701] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[1702] <= 32'b010010_11110_00001_1111111111111100; 	// sw
		disk[1703] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[1704] <= 32'b010010_11110_01111_1111111111111111; 	// sw
		disk[1705] <= 32'b010000_00000_10000_0000000000000001; 	// li
		disk[1706] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[1707] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[1708] <= 32'b010010_11110_10001_1111111111111101; 	// sw
		disk[1709] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[1710] <= 32'b001111_11110_00110_1111111111111100; 	// lw
		disk[1711] <= 32'b000000_00101_00110_10010_00000_001111; 	// let
		disk[1712] <= 32'b010101_10010_00000_0000000000100000; 	// jf
		disk[1713] <= 32'b010000_00000_10100_0000000000000001; 	// li
		disk[1714] <= 32'b000000_00101_10100_10011_00000_001111; 	// let
		disk[1715] <= 32'b010101_10011_00000_0000000000010010; 	// jf
		disk[1716] <= 32'b010010_11110_00101_1111111111111110; 	// sw
		disk[1717] <= 32'b111100_00000000000000000000011011; 	// j
		disk[1718] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1719] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[1720] <= 32'b000000_00101_00110_10101_00000_000000; 	// add
		disk[1721] <= 32'b010010_11110_10101_1111111111111110; 	// sw
		disk[1722] <= 32'b010010_11110_00110_1111111111111111; 	// sw
		disk[1723] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1724] <= 32'b001111_11110_00111_1111111111111110; 	// lw
		disk[1725] <= 32'b010010_11110_00111_0000000000000000; 	// sw
		disk[1726] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[1727] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[1728] <= 32'b000001_00101_10110_0000000000000001; 	// addi
		disk[1729] <= 32'b010010_11110_10110_1111111111111101; 	// sw
		disk[1730] <= 32'b001111_11110_00101_1111111111111101; 	// lw
		disk[1731] <= 32'b111100_00000000000000000000001001; 	// j
		disk[1732] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[1733] <= 32'b001110_00101_11001_0000000000000000; 	// mov
		disk[1734] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1735] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[1736] <= 32'b010000_00000_01111_0000000000001011; 	// li
		disk[1737] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[1738] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1739] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1740] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1741] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[1742] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[1743] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1744] <= 32'b001110_11001_00101_0000000000000000; 	// mov
		disk[1745] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1746] <= 32'b010000_00000_00010_0000000000000000; 	// li
		disk[1747] <= 32'b010100_00000_00001_0000000000000000; 	// out
		disk[1748] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[1749] <= 32'b011111_11111_00000_0000000000000000; 	// syscall
		
		// PROGRAMA 2
		disk[1800] <= 32'b111101_00000000000000000000100001;		// Jump to Main
		disk[1801] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[1802] <= 32'b010010_11110_00001_1111111111111100; 	// sw
		disk[1803] <= 32'b010010_11110_00010_1111111111111101; 	// sw
		disk[1804] <= 32'b010000_00000_01111_0000000000000000; 	// li
		disk[1805] <= 32'b010010_11110_01111_1111111111111110; 	// sw
		disk[1806] <= 32'b010000_00000_10000_0000000000000000; 	// li
		disk[1807] <= 32'b010010_11110_10000_0000000000000000; 	// sw
		disk[1808] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[1809] <= 32'b001111_11110_00110_1111111111111101; 	// lw
		disk[1810] <= 32'b000000_00101_00110_10001_00000_001110; 	// lt
		disk[1811] <= 32'b010101_10001_00000_0000000000011100; 	// jf
		disk[1812] <= 32'b001111_11110_00111_1111111111111100; 	// lw
		disk[1813] <= 32'b000000_00111_00101_10010_00000_000000; 	// add
		disk[1814] <= 32'b001111_10010_10010_0000000000000000; 	// lw
		disk[1815] <= 32'b001111_11110_01000_0000000000000000; 	// lw
		disk[1816] <= 32'b000000_01000_10010_10011_00000_001110; 	// lt
		disk[1817] <= 32'b010101_10011_00000_0000000000010111; 	// jf
		disk[1818] <= 32'b000000_00111_00101_10100_00000_000000; 	// add
		disk[1819] <= 32'b001111_10100_10100_0000000000000000; 	// lw
		disk[1820] <= 32'b010010_11110_10100_0000000000000000; 	// sw
		disk[1821] <= 32'b001111_11110_01000_0000000000000000; 	// lw
		disk[1822] <= 32'b010010_11110_00101_1111111111111111; 	// sw
		disk[1823] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[1824] <= 32'b000001_00101_10101_0000000000000001; 	// addi
		disk[1825] <= 32'b010010_11110_10101_1111111111111110; 	// sw
		disk[1826] <= 32'b001111_11110_00101_1111111111111110; 	// lw
		disk[1827] <= 32'b111100_00000000000000000000001000; 	// j
		disk[1828] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1829] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1830] <= 32'b010000_00000_00010_0000000000000001; 	// li
		disk[1831] <= 32'b010100_00000_00001_0000000000000001; 	// out
		disk[1832] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1833] <= 32'b000001_11110_11110_0000000000000111; 	// addi
		disk[1834] <= 32'b010001_11110_00101_1111111111111011; 	// la
		disk[1835] <= 32'b010000_00000_01111_0000000000001100; 	// li
		disk[1836] <= 32'b010010_00101_01111_0000000000000000; 	// sw
		disk[1837] <= 32'b010000_00000_10000_0000000000101001; 	// li
		disk[1838] <= 32'b010010_00101_10000_0000000000000001; 	// sw
		disk[1839] <= 32'b010000_00000_10001_0000000000010111; 	// li
		disk[1840] <= 32'b010010_00101_10001_0000000000000010; 	// sw
		disk[1841] <= 32'b010000_00000_10010_0000000001100010; 	// li
		disk[1842] <= 32'b010010_00101_10010_0000000000000011; 	// sw
		disk[1843] <= 32'b010000_00000_10011_0000000000100001; 	// li
		disk[1844] <= 32'b010010_00101_10011_0000000000000100; 	// sw
		disk[1845] <= 32'b010000_00000_10100_0000000000010101; 	// li
		disk[1846] <= 32'b010010_00101_10100_0000000000000101; 	// sw
		disk[1847] <= 32'b010001_11110_00001_1111111111111011; 	// la
		disk[1848] <= 32'b010000_00000_00010_0000000000000110; 	// li
		disk[1849] <= 32'b010010_11110_11111_1111111111111010; 	// sw
		disk[1850] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[1851] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[1852] <= 32'b001111_11110_11111_1111111111111010; 	// lw
		disk[1853] <= 32'b001110_11001_00101_0000000000000000; 	// mov
		disk[1854] <= 32'b000010_11110_11110_0000000000000111; 	// subi
		disk[1855] <= 32'b011111_11111_00000_0000000000000000; 	// syscall
		
		// PROGRAMA 3
		disk[1900] <= 32'b111101_00000000000000000000010100;		// Jump to Main
		disk[1901] <= 32'b000001_11110_11110_0000000000000100; 	// addi
		disk[1902] <= 32'b010010_11110_00001_1111111111111111; 	// sw
		disk[1903] <= 32'b010000_00000_01111_0000000000000001; 	// li
		disk[1904] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[1905] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1906] <= 32'b010000_00000_10001_0000000000000000; 	// li
		disk[1907] <= 32'b000000_00101_10001_10000_00000_010000; 	// gt
		disk[1908] <= 32'b010101_10000_00000_0000000000010001; 	// jf
		disk[1909] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[1910] <= 32'b000000_00110_00101_10010_00000_000010; 	// mul
		disk[1911] <= 32'b010010_11110_10010_0000000000000000; 	// sw
		disk[1912] <= 32'b001111_11110_00110_0000000000000000; 	// lw
		disk[1913] <= 32'b000010_00101_10011_0000000000000001; 	// subi
		disk[1914] <= 32'b010010_11110_10011_1111111111111111; 	// sw
		disk[1915] <= 32'b001111_11110_00101_1111111111111111; 	// lw
		disk[1916] <= 32'b111100_00000000000000000000000101; 	// j
		disk[1917] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1918] <= 32'b001110_00101_11001_0000000000000000; 	// mov
		disk[1919] <= 32'b000000_11111_00000_00000_00000_010010; 	// jr
		disk[1920] <= 32'b000001_11110_11110_0000000000000010; 	// addi
		disk[1921] <= 32'b010011_00000_01111_0000000000000000; 	// in
		disk[1922] <= 32'b010010_11110_01111_0000000000000000; 	// sw
		disk[1923] <= 32'b001111_11110_00101_0000000000000000; 	// lw
		disk[1924] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1925] <= 32'b010010_11110_11111_1111111111111111; 	// sw
		disk[1926] <= 32'b111110_00000000000000000000000001; 	// jal
		disk[1927] <= 32'b000010_11110_11110_0000000000000100; 	// subi
		disk[1928] <= 32'b001111_11110_11111_1111111111111111; 	// lw
		disk[1929] <= 32'b001110_11001_00101_0000000000000000; 	// mov
		disk[1930] <= 32'b001110_00101_00001_0000000000000000; 	// mov
		disk[1931] <= 32'b010000_00000_00010_0000000000000010; 	// li
		disk[1932] <= 32'b010100_00000_00001_0000000000000010; 	// out
		disk[1933] <= 32'b000010_11110_11110_0000000000000010; 	// subi
		disk[1934] <= 32'b011111_11111_00000_0000000000000000; 	// syscall

	end
endmodule
